----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
--
-- VHDL Architecture conv_lib.conv_mult.scm
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 17:37:47 26/04/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library dsp_prim_lib;

library conv_lib;

architecture scm of conv_mult is

  -- Architecture declarations

  -- Internal signal declarations
  signal CLKEN  : std_logic;                       -- ena
  signal IDATA1 : std_logic_vector(31 downto 0);
  signal RDATA1 : std_logic_vector(31 downto 0);   -- az
  signal RST    : std_logic;                       -- aclr
  signal SYNC   : std_logic;


  -- Component Declarations
  component retime
  generic (
    dataw_g  : natural;
    stages_g : natural
  );
  port (
    DATA    : in     std_logic_vector (dataw_g-1 downto 0);
    DE      : in     std_logic ;
    SYNC    : in     std_logic ;
    CLK     : in     std_logic ;
    CLKEN   : in     std_logic ;
    RST_N   : in     std_logic ;
    DATAOUT : out    std_logic_vector (dataw_g-1 downto 0);
    DEOUT   : out    std_logic 
  );
  end component retime;
  component cmplxmult_fp
  port (
    ACLR        : in     std_logic ;                     -- aclr
    AY_IM       : in     std_logic_vector (31 downto 0); -- ax
    AY_RE       : in     std_logic_vector (31 downto 0); -- ax
    AZ_IM       : in     std_logic_vector (31 downto 0); -- az
    AZ_RE       : in     std_logic_vector (31 downto 0); -- az
    CLK         : in     std_logic ;                     -- clk
    ENA         : in     std_logic ;                     -- ena
    CHAINOUT_IM : out    std_logic_vector (31 downto 0); -- result
    CHAINOUT_RE : out    std_logic_vector (31 downto 0); -- result
    RESULT_IM   : out    std_logic_vector (31 downto 0); -- result
    RESULT_RE   : out    std_logic_vector (31 downto 0)  -- result
  );
  end component cmplxmult_fp;

  -- Optional embedded configurations
  -- pragma synthesis_off
  for all : cmplxmult_fp use entity dsp_prim_lib.cmplxmult_fp;
  for all : retime use entity conv_lib.retime;
  -- pragma synthesis_on


begin
  -- Architecture concurrent statements
  -- HDL Embedded Text Block 1 eb1
  -- eb1 1
  CLKEN <= '1';
  RST <= not RST_SYS_N;
  SYNC <= '0';                                  


  -- Instance port mappings.
  idatain_i : retime
    generic map (
      dataw_g  => 32,
      stages_g => 1
    )
    port map (
      DATA    => IDATA,
      DE      => VALID,
      SYNC    => SYNC,
      CLK     => CLK_SYS,
      CLKEN   => CLKEN,
      RST_N   => RST_SYS_N,
      DATAOUT => IDATA1,
      DEOUT   => open
    );
  rdatain_i : retime
    generic map (
      dataw_g  => 32,
      stages_g => 1
    )
    port map (
      DATA    => RDATA,
      DE      => VALID,
      SYNC    => SYNC,
      CLK     => CLK_SYS,
      CLKEN   => CLKEN,
      RST_N   => RST_SYS_N,
      DATAOUT => RDATA1,
      DEOUT   => open
    );
  --  Module Name:  CMPLXMULT
  --
  --  Source Path:  cmplxmult.vhd
  --
  --  Description:
  --
  --  Author:       jon.taylor@covnetics.com
  --
  -- --------------------------------------------------------------------------
  --  Rev  Auth     Date      Revision History
  --
  --  0.1  JT     26/11/2015  Initial revision.
  -- --------------------------------------------------------------------------
  --        __
  --     ,/'__`\                             _     _
  --    ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
  --    ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
  --    '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
  --     '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
  --
  --  Copyright (c) Covnetics Limited 2015 All Rights Reserved. The information
  --  contained herein remains the property of Covnetics Limited and may not be
  --  copied or reproduced in any format or medium without the written consent
  --  of Covnetics Limited.
  --
  -- --------------------------------------------------------------------------
  --  VHDL Version: VHDL '93
  -- --------------------------------------------------------------------------
  --
  --  Module Name:  CMPLXMULT
  -- 
  --  Source Path:  cmplxmult.vhd
  -- 
  --  Description:  
  -- 
  --  Author:       jon.taylor@covnetics.com
  -- 
  -- --------------------------------------------------------------------------
  --  Rev  Auth     Date      Revision History
  -- 
  --  0.1  JT     26/11/2015  Initial revision.
  -- --------------------------------------------------------------------------
  --        __
  --     ,/'__`\                             _     _
  --    ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
  --    ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
  --    '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
  --     '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
  -- 
  --  Copyright (c) Covnetics Limited 2015 All Rights Reserved. The information
  --  contained herein remains the property of Covnetics Limited and may not be
  --  copied or reproduced in any format or medium without the written consent
  --  of Covnetics Limited.
  -- 
  -- --------------------------------------------------------------------------
  --  VHDL Version: VHDL '93
  -- --------------------------------------------------------------------------
  -- 
  cmplx_mult_conj_i : cmplxmult_fp
    port map (
      ACLR        => RST,
      AY_IM       => ICOEFCONJ,
      AY_RE       => RCOEFCONJ,
      AZ_IM       => IDATA1,
      AZ_RE       => RDATA1,
      CLK         => CLK_SYS,
      ENA         => CLKEN,
      CHAINOUT_IM => open,
      CHAINOUT_RE => open,
      RESULT_IM   => IDATACONJOUT,
      RESULT_RE   => RDATACONJOUT
    );
  --  Module Name:  CMPLXMULT
  --
  --  Source Path:  cmplxmult.vhd
  --
  --  Description:
  --
  --  Author:       jon.taylor@covnetics.com
  --
  -- --------------------------------------------------------------------------
  --  Rev  Auth     Date      Revision History
  --
  --  0.1  JT     26/11/2015  Initial revision.
  -- --------------------------------------------------------------------------
  --        __
  --     ,/'__`\                             _     _
  --    ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
  --    ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
  --    '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
  --     '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
  --
  --  Copyright (c) Covnetics Limited 2015 All Rights Reserved. The information
  --  contained herein remains the property of Covnetics Limited and may not be
  --  copied or reproduced in any format or medium without the written consent
  --  of Covnetics Limited.
  --
  -- --------------------------------------------------------------------------
  --  VHDL Version: VHDL '93
  -- --------------------------------------------------------------------------
  --
  --  Module Name:  CMPLXMULT
  -- 
  --  Source Path:  cmplxmult.vhd
  -- 
  --  Description:  
  -- 
  --  Author:       jon.taylor@covnetics.com
  -- 
  -- --------------------------------------------------------------------------
  --  Rev  Auth     Date      Revision History
  -- 
  --  0.1  JT     26/11/2015  Initial revision.
  -- --------------------------------------------------------------------------
  --        __
  --     ,/'__`\                             _     _
  --    ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
  --    ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
  --    '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
  --     '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
  -- 
  --  Copyright (c) Covnetics Limited 2015 All Rights Reserved. The information
  --  contained herein remains the property of Covnetics Limited and may not be
  --  copied or reproduced in any format or medium without the written consent
  --  of Covnetics Limited.
  -- 
  -- --------------------------------------------------------------------------
  --  VHDL Version: VHDL '93
  -- --------------------------------------------------------------------------
  -- 
  cmplx_mult_i : cmplxmult_fp
    port map (
      ACLR        => RST,
      AY_IM       => ICOEF,
      AY_RE       => RCOEF,
      AZ_IM       => IDATA1,
      AZ_RE       => RDATA1,
      CLK         => CLK_SYS,
      ENA         => CLKEN,
      CHAINOUT_IM => open,
      CHAINOUT_RE => open,
      RESULT_IM   => IDATAOUT,
      RESULT_RE   => RDATAOUT
    );

end architecture scm;
