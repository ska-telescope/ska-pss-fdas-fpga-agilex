-- mult_fp_co.vhd

-- Generated using ACDS version 22.2 94

library IEEE;
library s20_native_floating_point_dsp_1910;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mult_fp_co is
	port (
		fp32_mult_a   : in  std_logic_vector(31 downto 0) := (others => '0'); --   fp32_mult_a.fp32_mult_a
		fp32_mult_b   : in  std_logic_vector(31 downto 0) := (others => '0'); --   fp32_mult_b.fp32_mult_b
		clr0          : in  std_logic                     := '0';             --          clr0.reset
		clr1          : in  std_logic                     := '0';             --          clr1.reset
		clk           : in  std_logic                     := '0';             --           clk.clk
		ena           : in  std_logic_vector(2 downto 0)  := (others => '0'); --           ena.ena
		fp32_result   : out std_logic_vector(31 downto 0);                    --   fp32_result.fp32_result
		fp32_chainout : out std_logic_vector(31 downto 0)                     -- fp32_chainout.fp32_chainout
	);
end entity mult_fp_co;

architecture rtl of mult_fp_co is
	component mult_fp_co_s20_native_floating_point_dsp_1910_nhmydci_cmp is
		port (
			fp32_mult_a   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- fp32_mult_a
			fp32_mult_b   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- fp32_mult_b
			clr0          : in  std_logic                     := 'X';             -- reset
			clr1          : in  std_logic                     := 'X';             -- reset
			clk           : in  std_logic                     := 'X';             -- clk
			ena           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- ena
			fp32_result   : out std_logic_vector(31 downto 0);                    -- fp32_result
			fp32_chainout : out std_logic_vector(31 downto 0)                     -- fp32_chainout
		);
	end component mult_fp_co_s20_native_floating_point_dsp_1910_nhmydci_cmp;

	for s20_native_floating_point_dsp_0 : mult_fp_co_s20_native_floating_point_dsp_1910_nhmydci_cmp
		use entity s20_native_floating_point_dsp_1910.mult_fp_co_s20_native_floating_point_dsp_1910_nhmydci;
begin

	s20_native_floating_point_dsp_0 : component mult_fp_co_s20_native_floating_point_dsp_1910_nhmydci_cmp
		port map (
			fp32_mult_a   => fp32_mult_a,   --   fp32_mult_a.fp32_mult_a
			fp32_mult_b   => fp32_mult_b,   --   fp32_mult_b.fp32_mult_b
			clr0          => clr0,          --          clr0.reset
			clr1          => clr1,          --          clr1.reset
			clk           => clk,           --           clk.clk
			ena           => ena,           --           ena.ena
			fp32_result   => fp32_result,   --   fp32_result.fp32_result
			fp32_chainout => fp32_chainout  -- fp32_chainout.fp32_chainout
		);

end architecture rtl; -- of mult_fp_co
