----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity cld_lib.dual_port_ram.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 13:26:50 13/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library cld_lib;
use cld_lib.all;

ENTITY dual_port_ram IS
  GENERIC( 
    abits_g : integer;
    dbits_g : integer
  );
  PORT( 
    aa    : IN     std_logic_vector (abits_g-1 DOWNTO 0);
    ai    : IN     std_logic_vector (dbits_g-1 DOWNTO 0);
    awren : IN     std_logic;
    ba    : IN     std_logic_vector (abits_g-1 DOWNTO 0);
    clk   : IN     std_logic;
    bo    : OUT    std_logic_vector (dbits_g-1 DOWNTO 0)
  );

-- Declarations

END ENTITY dual_port_ram ;

