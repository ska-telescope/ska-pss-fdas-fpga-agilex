----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.conv_ifft_ctrl.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 19:09:50 11/07/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity conv_ifft_ctrl is
  generic( 
    stages_g    : natural;
    loop_g      : natural;    --lte 2**loop_bits_g
    loop_bits_g : natural
  );
  port( 
    SOF          : in     std_logic;
    EOF          : in     std_logic;
    VALID        : in     std_logic;
    READY        : in     std_logic;
    SYNC         : in     std_logic;
    LOOP_NUM     : in     std_logic_vector (loop_bits_g downto 0);
    CLK          : in     std_logic;
    CLKEN        : in     std_logic;
    RST_N        : in     std_logic;
    SOFOUT       : out    std_logic;
    EOFOUT       : out    std_logic;
    VALIDOUT     : out    std_logic;
    LOOP_ADDROUT : out    std_logic_vector (loop_bits_g-1 downto 0);
    WRENOUT      : out    std_logic_vector (loop_g-1 downto 0)
  );

-- Declarations

end entity conv_ifft_ctrl ;

