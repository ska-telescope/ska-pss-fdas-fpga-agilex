----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
--
-- VHDL Architecture cld_lib.cld.scm
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 13:26:51 13/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library cld_lib;
use cld_lib.all;


ARCHITECTURE scm OF cld IS

  -- Architecture declarations

  -- Internal signal declarations
  SIGNAL completed_read_sample_s : std_logic_vector(sample_count_width_g -1 DOWNTO 0);
  SIGNAL ddr_done_s              : std_logic;
  SIGNAL ddr_en_s                : std_logic;
  SIGNAL ddr_reading_finished_s  : std_logic;
  SIGNAL fft_zeros_s             : std_logic;
  SIGNAL fifo_raddr_s            : std_logic_vector(fifo_raddr_width_g -1  DOWNTO 0);
  SIGNAL fifo_waddr_s            : std_logic_vector(fifo_waddr_width_g -1  DOWNTO 0);
  SIGNAL wait_req_s              : std_logic;
  SIGNAL write_sample_s          : std_logic_vector(sample_count_width_g -1 DOWNTO 0);


  -- Component Declarations
  COMPONENT cld_ddr_rag
  GENERIC (
    fft_ddr_addr_num_g       : integer;
    fft_ddr_addr_num_width_g : integer;
    fop_ddr_addr_max_width_g : integer
  );
  PORT (
    cld_enable   : IN     std_logic ;
    cld_page     : IN     std_logic_vector (31 DOWNTO 0);
    cld_trigger  : IN     std_logic ;
    clk_sys      : IN     std_logic ;
    data_valid   : IN     std_logic ;
    ddr_en       : IN     std_logic ;
    rst_sys_n    : IN     std_logic ;
    wait_request : IN     std_logic ;
    ddr_addr     : OUT    std_logic_vector (31 DOWNTO 0);
    ddr_done     : OUT    std_logic ;
    ddr_read     : OUT    std_logic 
  );
  END COMPONENT cld_ddr_rag;
  COMPONENT cld_fifo
  GENERIC (
    fifo_waddr_width_g : integer;
    fifo_raddr_width_g : integer;
    ddr_g              : integer
  );
  PORT (
    clk_sys      : IN     std_logic ;
    data_valid   : IN     std_logic ;
    ddr_data     : IN     std_logic_vector (512*ddr_g -1  DOWNTO 0);
    fft_zeros    : IN     std_logic ;
    fifo_raddr_s : IN     std_logic_vector (fifo_raddr_width_g -1  DOWNTO 0);
    fifo_waddr_s : IN     std_logic_vector (fifo_waddr_width_g -1  DOWNTO 0);
    rst_sys_n    : IN     std_logic ;
    wait_req     : IN     std_logic ;
    conv_data    : OUT    std_logic_vector (63  DOWNTO 0)
  );
  END COMPONENT cld_fifo;
  COMPONENT cld_fifo_rag
  GENERIC (
    fifo_raddr_width_g   : integer;
    fft_count_width_g    : integer;
    sample_count_width_g : integer;
    fft_g                : integer;
    ddr_g                : integer
  );
  PORT (
    cld_enable            : IN     std_logic ;
    cld_trigger           : IN     std_logic ;
    clk_sys               : IN     std_logic ;
    ddr_reading_finished  : IN     std_logic ;
    fop_sample_num        : IN     std_logic_vector (22 DOWNTO 0);
    overlap_int           : IN     std_logic_vector (4 DOWNTO 0);
    overlap_rem           : IN     std_logic_vector (4 DOWNTO 0);
    overlap_size          : IN     std_logic_vector (9  DOWNTO 0);
    ready                 : IN     std_logic ;
    rst_sys_n             : IN     std_logic ;
    write_sample          : IN     std_logic_vector (sample_count_width_g -1 DOWNTO 0);
    cld_done              : OUT    std_logic ;
    completed_read_sample : OUT    std_logic_vector (sample_count_width_g -1 DOWNTO 0);
    conv_req              : OUT    std_logic ;
    eof                   : OUT    std_logic ;
    fft_sample            : OUT    std_logic_vector (fft_count_width_g-1  DOWNTO 0);
    fft_zeros             : OUT    std_logic ;
    fifo_raddr            : OUT    std_logic_vector (fifo_raddr_width_g -1  DOWNTO 0);
    sof                   : OUT    std_logic ;
    valid                 : OUT    std_logic ;
    wait_req              : OUT    std_logic 
  );
  END COMPONENT cld_fifo_rag;
  COMPONENT cld_fifo_wag
  GENERIC (
    fifo_waddr_width_g   : integer;
    fft_count_width_g    : integer;
    sample_count_width_g : integer;
    fft_g                : integer;
    ddr_g                : integer
  );
  PORT (
    cld_enable            : IN     std_logic ;
    cld_trigger           : IN     std_logic ;
    clk_sys               : IN     std_logic ;
    completed_read_sample : IN     std_logic_vector (sample_count_width_g -1 DOWNTO 0);
    data_valid            : IN     std_logic ;
    ddr_done              : IN     std_logic ;
    fop_sample_num        : IN     std_logic_vector (22 DOWNTO 0);
    rst_sys_n             : IN     std_logic ;
    ddr_en                : OUT    std_logic ;
    ddr_reading_finished  : OUT    std_logic ;
    fifo_waddr            : OUT    std_logic_vector (fifo_waddr_width_g -1  DOWNTO 0);
    write_sample          : OUT    std_logic_vector (sample_count_width_g -1 DOWNTO 0)
  );
  END COMPONENT cld_fifo_wag;

  -- Optional embedded configurations
  -- pragma synthesis_off
  FOR ALL : cld_ddr_rag USE ENTITY cld_lib.cld_ddr_rag;
  FOR ALL : cld_fifo USE ENTITY cld_lib.cld_fifo;
  FOR ALL : cld_fifo_rag USE ENTITY cld_lib.cld_fifo_rag;
  FOR ALL : cld_fifo_wag USE ENTITY cld_lib.cld_fifo_wag;
  -- pragma synthesis_on


BEGIN

  -- Instance port mappings.
  cld_ddr_rag_1 : cld_ddr_rag
    GENERIC MAP (
      fft_ddr_addr_num_g       => fft_ddr_addr_num_g,
      fft_ddr_addr_num_width_g => fft_ddr_addr_num_width_g,
      fop_ddr_addr_max_width_g => fop_ddr_addr_max_width_g
    )
    PORT MAP (
      cld_enable   => cld_enable,
      cld_page     => cld_page,
      cld_trigger  => cld_trigger,
      clk_sys      => clk_sys,
      data_valid   => data_valid,
      ddr_en       => ddr_en_s,
      rst_sys_n    => rst_sys_n,
      wait_request => wait_request,
      ddr_addr     => ddr_addr,
      ddr_done     => ddr_done_s,
      ddr_read     => ddr_read
    );
  cld_fifo_1 : cld_fifo
    GENERIC MAP (
      fifo_waddr_width_g => fifo_waddr_width_g,
      fifo_raddr_width_g => fifo_raddr_width_g,
      ddr_g              => ddr_g
    )
    PORT MAP (
      clk_sys      => clk_sys,
      data_valid   => data_valid,
      ddr_data     => ddr_data,
      fft_zeros    => fft_zeros_s,
      fifo_raddr_s => fifo_raddr_s,
      fifo_waddr_s => fifo_waddr_s,
      rst_sys_n    => rst_sys_n,
      wait_req     => wait_req_s,
      conv_data    => conv_data
    );
  cld_fifo_rag_1 : cld_fifo_rag
    GENERIC MAP (
      fifo_raddr_width_g   => fifo_raddr_width_g,
      fft_count_width_g    => fft_count_width_g,
      sample_count_width_g => sample_count_width_g,
      fft_g                => fft_g,
      ddr_g                => ddr_g
    )
    PORT MAP (
      cld_enable            => cld_enable,
      cld_trigger           => cld_trigger,
      clk_sys               => clk_sys,
      ddr_reading_finished  => ddr_reading_finished_s,
      fop_sample_num        => fop_sample_num,
      overlap_int           => overlap_int,
      overlap_rem           => overlap_rem,
      overlap_size          => overlap_size,
      ready                 => ready,
      rst_sys_n             => rst_sys_n,
      write_sample          => write_sample_s,
      cld_done              => cld_done,
      completed_read_sample => completed_read_sample_s,
      conv_req              => conv_req,
      eof                   => eof,
      fft_sample            => fft_sample,
      fft_zeros             => fft_zeros_s,
      fifo_raddr            => fifo_raddr_s,
      sof                   => sof,
      valid                 => valid,
      wait_req              => wait_req_s
    );
  cld_fifo_wag_1 : cld_fifo_wag
    GENERIC MAP (
      fifo_waddr_width_g   => fifo_waddr_width_g,
      fft_count_width_g    => fft_count_width_g,
      sample_count_width_g => sample_count_width_g,
      fft_g                => fft_g,
      ddr_g                => ddr_g
    )
    PORT MAP (
      cld_enable            => cld_enable,
      cld_trigger           => cld_trigger,
      clk_sys               => clk_sys,
      completed_read_sample => completed_read_sample_s,
      data_valid            => data_valid,
      ddr_done              => ddr_done_s,
      fop_sample_num        => fop_sample_num,
      rst_sys_n             => rst_sys_n,
      ddr_en                => ddr_en_s,
      ddr_reading_finished  => ddr_reading_finished_s,
      fifo_waddr            => fifo_waddr_s,
      write_sample          => write_sample_s
    );

END ARCHITECTURE scm;
