----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.conv_result_str.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 11:05:59 13/05/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity conv_result_str is
  generic( 
    dbits_g  : natural;
    depth_g  : natural;
    abits_g  : natural;
    pages_g  : natural;    -- lte 2**(pgbits_g-1)
    pgbits_g : natural
  );
  port( 
    CLK_SYS   : in     std_logic;
    RST_SYS_N : in     std_logic;
    RDADDR    : in     std_logic_vector (abits_g-1 downto 0);
    RDEN      : in     std_logic;
    RDEOF     : in     std_logic;
    DATAOUT   : out    std_logic_vector (dbits_g-1 downto 0);
    DATA      : in     std_logic_vector (dbits_g-1 downto 0);
    VALID     : in     std_logic;
    SOF       : in     std_logic;
    EOF       : in     std_logic;
    SYNC      : in     std_logic;
    AVAILOUT  : out    std_logic;
    READYOUT  : out    std_logic;
    OVERFLOW  : out    std_logic;
    DONEOUT   : out    std_logic
  );

-- Declarations

end entity conv_result_str ;

