----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
--
-- VHDL Architecture conv_lib.conv_pwr.scm
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 09:38:51 11/05/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library conv_lib;
library dsp_prim_lib;

architecture scm of conv_pwr is

  -- Architecture declarations

  -- Internal signal declarations
  signal ACLR     : std_logic;                       -- aclr
  signal CLKEN    : std_logic_vector(2 downto 0);
  signal CTRL     : std_logic_vector(1 downto 0);
  signal CTRLOUT  : std_logic_vector(1 downto 0);
  signal RTCLKEN  : std_logic;
  signal chainout : std_logic_vector(31 downto 0);   -- chainout.chainout


  -- Component Declarations
  component retime
  generic (
    dataw_g  : natural;
    stages_g : natural
  );
  port (
    DATA    : in     std_logic_vector (dataw_g-1 downto 0);
    DE      : in     std_logic ;
    SYNC    : in     std_logic ;
    CLK     : in     std_logic ;
    CLKEN   : in     std_logic ;
    RST_N   : in     std_logic ;
    DATAOUT : out    std_logic_vector (dataw_g-1 downto 0);
    DEOUT   : out    std_logic 
  );
  end component retime;
  component mult_fp_co
  port (
    clr0          : in     std_logic                      := '0';
    fp32_mult_a   : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_mult_b   : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_chainout : out    std_logic_vector (31 downto 0);
    clk           : in     std_logic                      := '0';
    ena           : in     std_logic_vector (2 downto 0)  := (others => '0');
    fp32_result   : out    std_logic_vector (31 downto 0);
    clr1          : in     std_logic                      := '0'
  );
  end component mult_fp_co;
  component multadd_fp_ci
  port (
    clr0         : in     std_logic                      := '0';
    fp32_mult_a  : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_mult_b  : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_chainin : in     std_logic_vector (31 downto 0) := (others => '0');
    clk          : in     std_logic                      := '0';
    ena          : in     std_logic_vector (2 downto 0)  := (others => '0');
    fp32_result  : out    std_logic_vector (31 downto 0);
    clr1         : in     std_logic                      := '0'
  );
  end component multadd_fp_ci;

  -- Optional embedded configurations
  -- pragma synthesis_off
  for all : mult_fp_co use entity dsp_prim_lib.mult_fp_co;
  for all : multadd_fp_ci use entity dsp_prim_lib.multadd_fp_ci;
  for all : retime use entity conv_lib.retime;
  -- pragma synthesis_on


begin
  -- Architecture concurrent statements
  -- HDL Embedded Text Block 1 eb1
  -- eb1 1
  CLKEN <= (others => '1');
  RTCLKEN <= '1';
  ACLR <= not RST_SYS_N;
  CTRL <= EOF & SOF;
  SOFOUT <= CTRLOUT(0);
  EOFOUT <= CTRLOUT(1);


  -- Instance port mappings.
  retime_i : retime
    generic map (
      dataw_g  => 2,
      stages_g => 4
    )
    port map (
      DATA    => CTRL,
      DE      => VALID,
      SYNC    => SYNC,
      CLK     => CLK_SYS,
      CLKEN   => RTCLKEN,
      RST_N   => RST_SYS_N,
      DATAOUT => CTRLOUT,
      DEOUT   => VALIDOUT
    );
  mult_i : mult_fp_co
    port map (
      clr0          => ACLR,
      fp32_mult_a   => RDATA,
      fp32_mult_b   => RDATA,
      fp32_chainout => chainout,
      clk           => CLK_SYS,
      ena           => CLKEN,
      fp32_result   => open,
      clr1          => ACLR
    );
  multadd_i : multadd_fp_ci
    port map (
      clr0         => ACLR,
      fp32_mult_a  => IDATA,
      fp32_mult_b  => IDATA,
      fp32_chainin => chainout,
      clk          => CLK_SYS,
      ena          => CLKEN,
      fp32_result  => DATAOUT,
      clr1         => ACLR
    );

end architecture scm;
