----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.conv_pwr.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 17:39:18 26/04/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity conv_pwr is
  port( 
    CLK_SYS   : in     std_logic;
    EOF       : in     std_logic;
    IDATA     : in     std_logic_vector (31 downto 0);  -- az
    RDATA     : in     std_logic_vector (31 downto 0);
    RST_SYS_N : in     std_logic;
    SOF       : in     std_logic;
    SYNC      : in     std_logic;
    VALID     : in     std_logic;
    DATAOUT   : out    std_logic_vector (31 downto 0);
    EOFOUT    : out    std_logic;
    SOFOUT    : out    std_logic;
    VALIDOUT  : out    std_logic
  );

-- Declarations

end entity conv_pwr ;

