module RESET_RELEASE (
		output wire  ninit_done  // ninit_done.ninit_done
	);
endmodule

