----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity cld_lib.cld_fifo.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 13:26:50 13/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY cld_fifo IS
  GENERIC( 
    fifo_waddr_width_g : integer;
    fifo_raddr_width_g : integer;
    ddr_g              : integer
  );
  PORT( 
    clk_sys      : IN     std_logic;
    data_valid   : IN     std_logic;
    ddr_data     : IN     std_logic_vector (512*ddr_g -1  DOWNTO 0);
    fft_zeros    : IN     std_logic;
    fifo_raddr_s : IN     std_logic_vector (fifo_raddr_width_g -1  DOWNTO 0);
    fifo_waddr_s : IN     std_logic_vector (fifo_waddr_width_g -1  DOWNTO 0);
    rst_sys_n    : IN     std_logic;
    wait_req     : IN     std_logic;
    conv_data    : OUT    std_logic_vector (63  DOWNTO 0)
  );

-- Declarations

END ENTITY cld_fifo ;

