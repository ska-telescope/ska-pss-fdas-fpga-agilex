-- multsub_fp_ci.vhd

-- Generated using ACDS version 22.2 94

library IEEE;
library s20_native_floating_point_dsp_1910;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity multsub_fp_ci is
	port (
		fp32_mult_a  : in  std_logic_vector(31 downto 0) := (others => '0'); --  fp32_mult_a.fp32_mult_a
		fp32_mult_b  : in  std_logic_vector(31 downto 0) := (others => '0'); --  fp32_mult_b.fp32_mult_b
		fp32_chainin : in  std_logic_vector(31 downto 0) := (others => '0'); -- fp32_chainin.fp32_chainin
		clr0         : in  std_logic                     := '0';             --         clr0.reset
		clr1         : in  std_logic                     := '0';             --         clr1.reset
		clk          : in  std_logic                     := '0';             --          clk.clk
		ena          : in  std_logic_vector(2 downto 0)  := (others => '0'); --          ena.ena
		fp32_result  : out std_logic_vector(31 downto 0)                     --  fp32_result.fp32_result
	);
end entity multsub_fp_ci;

architecture rtl of multsub_fp_ci is
	component multsub_fp_ci_s20_native_floating_point_dsp_1910_xbnuxwa_cmp is
		port (
			fp32_mult_a  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- fp32_mult_a
			fp32_mult_b  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- fp32_mult_b
			fp32_chainin : in  std_logic_vector(31 downto 0) := (others => 'X'); -- fp32_chainin
			clr0         : in  std_logic                     := 'X';             -- reset
			clr1         : in  std_logic                     := 'X';             -- reset
			clk          : in  std_logic                     := 'X';             -- clk
			ena          : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- ena
			fp32_result  : out std_logic_vector(31 downto 0)                     -- fp32_result
		);
	end component multsub_fp_ci_s20_native_floating_point_dsp_1910_xbnuxwa_cmp;

	for s20_native_floating_point_dsp_0 : multsub_fp_ci_s20_native_floating_point_dsp_1910_xbnuxwa_cmp
		use entity s20_native_floating_point_dsp_1910.multsub_fp_ci_s20_native_floating_point_dsp_1910_xbnuxwa;
begin

	s20_native_floating_point_dsp_0 : component multsub_fp_ci_s20_native_floating_point_dsp_1910_xbnuxwa_cmp
		port map (
			fp32_mult_a  => fp32_mult_a,  --  fp32_mult_a.fp32_mult_a
			fp32_mult_b  => fp32_mult_b,  --  fp32_mult_b.fp32_mult_b
			fp32_chainin => fp32_chainin, -- fp32_chainin.fp32_chainin
			clr0         => clr0,         --         clr0.reset
			clr1         => clr1,         --         clr1.reset
			clk          => clk,          --          clk.clk
			ena          => ena,          --          ena.ena
			fp32_result  => fp32_result   --  fp32_result.fp32_result
		);

end architecture rtl; -- of multsub_fp_ci
