----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
--
-- VHDL Architecture dsp_prim_lib.cmplxmult_fp.scm
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 15:34:19 10/05/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;

library dsp_prim_lib;

architecture scm of cmplxmult_fp is

  -- Architecture declarations

  -- Internal signal declarations
  signal chainout  : std_logic_vector(31 downto 0);   -- chainout.chainout
  signal chainout1 : std_logic_vector(31 downto 0);   -- chainout.chainout
  signal ena_s     : std_logic_vector(2 downto 0);


  -- Component Declarations
  component mult_fp_co
  port (
    clr0          : in     std_logic                      := '0';
    fp32_mult_a   : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_mult_b   : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_chainout : out    std_logic_vector (31 downto 0);
    clk           : in     std_logic                      := '0';
    ena           : in     std_logic_vector (2 downto 0)  := (others => '0');
    fp32_result   : out    std_logic_vector (31 downto 0);
    clr1          : in     std_logic                      := '0'
  );
  end component mult_fp_co;
  component multadd_fp_ci
  port (
    clr0         : in     std_logic                      := '0';
    fp32_mult_a  : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_mult_b  : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_chainin : in     std_logic_vector (31 downto 0) := (others => '0');
    clk          : in     std_logic                      := '0';
    ena          : in     std_logic_vector (2 downto 0)  := (others => '0');
    fp32_result  : out    std_logic_vector (31 downto 0);
    clr1         : in     std_logic                      := '0'
  );
  end component multadd_fp_ci;
  component multsub_fp_ci
  port (
    clr0         : in     std_logic                      := '0';
    fp32_mult_a  : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_mult_b  : in     std_logic_vector (31 downto 0) := (others => '0');
    fp32_chainin : in     std_logic_vector (31 downto 0) := (others => '0');
    clk          : in     std_logic                      := '0';
    ena          : in     std_logic_vector (2 downto 0)  := (others => '0');
    fp32_result  : out    std_logic_vector (31 downto 0);
    clr1         : in     std_logic                      := '0'
  );
  end component multsub_fp_ci;

  -- Optional embedded configurations
  -- pragma synthesis_off
  for all : mult_fp_co use entity dsp_prim_lib.mult_fp_co;
  for all : multadd_fp_ci use entity dsp_prim_lib.multadd_fp_ci;
  for all : multsub_fp_ci use entity dsp_prim_lib.multsub_fp_ci;
  -- pragma synthesis_on


begin
  -- Architecture concurrent statements
  -- HDL Embedded Text Block 1 eb1
  -- eb1 1 
  ena_s <= (others => ENA);                                      


  -- Instance port mappings.
  U_0 : mult_fp_co
    port map (
      clr0          => ACLR,
      fp32_mult_a   => AY_RE,
      fp32_mult_b   => AZ_IM,
      fp32_chainout => chainout,
      clk           => CLK,
      ena           => ena_s,
      fp32_result   => open,
      clr1          => ACLR
    );
  U_3 : mult_fp_co
    port map (
      clr0          => ACLR,
      fp32_mult_a   => AY_IM,
      fp32_mult_b   => AZ_IM,
      fp32_chainout => chainout1,
      clk           => CLK,
      ena           => ena_s,
      fp32_result   => open,
      clr1          => ACLR
    );
  U_1 : multadd_fp_ci
    port map (
      clr0         => ACLR,
      fp32_mult_a  => AY_IM,
      fp32_mult_b  => AZ_RE,
      fp32_chainin => chainout,
      clk          => CLK,
      ena          => ena_s,
      fp32_result  => RESULT_IM,
      clr1         => ACLR
    );
  U_2 : multsub_fp_ci
    port map (
      clr0         => ACLR,
      fp32_mult_a  => AY_RE,
      fp32_mult_b  => AZ_RE,
      fp32_chainin => chainout1,
      clk          => CLK,
      ena          => ena_s,
      fp32_result  => RESULT_RE,
      clr1         => ACLR
    );

end architecture scm;
