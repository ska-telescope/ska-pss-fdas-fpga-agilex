----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity cld_lib.cld_ddr_rag.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 13:26:50 13/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY cld_ddr_rag IS
  GENERIC( 
    fft_ddr_addr_num_g       : integer;
    fft_ddr_addr_num_width_g : integer;
    fop_ddr_addr_max_width_g : integer
  );
  PORT( 
    cld_enable   : IN     std_logic;
    cld_page     : IN     std_logic_vector (31 DOWNTO 0);
    cld_trigger  : IN     std_logic;
    clk_sys      : IN     std_logic;
    data_valid   : IN     std_logic;
    ddr_en       : IN     std_logic;
    rst_sys_n    : IN     std_logic;
    wait_request : IN     std_logic;
    ddr_addr     : OUT    std_logic_vector (31 DOWNTO 0);
    ddr_done     : OUT    std_logic;
    ddr_read     : OUT    std_logic
  );

-- Declarations

END ENTITY cld_ddr_rag ;

