----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.fop_str.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 19:00:22 11/07/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fop_str is
  generic( 
    ddr_g            : natural;
    abits_g          : natural;
    ifft_g           : natural;
    ifft_loop_g      : natural;    -- number of output frame repeats lte 2**ifft_loop_bits_g
    ifft_loop_bits_g : natural;
    fop_num_bits_g   : natural;
    delay_g          : natural;
    delaybits_g      : natural
  );
  port( 
    CLK_SYS       : in     std_logic;
    RST_SYS_N     : in     std_logic;
    RDADDROUT     : out    std_logic_vector (abits_g-1 downto 0);
    RDADDR0OUT    : out    std_logic_vector (abits_g-1 downto 0);
    RDENOUT       : out    std_logic_vector (2*ifft_g*ifft_loop_g downto 0);
    RDEOFOUT      : out    std_logic;
    RDDATA        : in     std_logic_vector ((2*ifft_g*ifft_loop_g+1)*32-1 downto 0);
    DDR_WAITREQ   : in     std_logic;
    AVAIL         : in     std_logic;
    DDR_ADDROUT   : out    std_logic_vector (25 downto 0);
    DDR_DATAOUT   : out    std_logic_vector (ddr_g*512-1 downto 0);
    DDR_VALIDOUT  : out    std_logic;
    DONEOUT       : out    std_logic;
    CONV_DONEOUT  : out    std_logic;
    IFFT_LOOP_NUM : in     std_logic_vector (ifft_loop_bits_g downto 0);
    FOP_NUM       : in     std_logic_vector (fop_num_bits_g-1 downto 0);
    OVERLAP_SIZE  : in     std_logic_vector (abits_g-1 downto 0);
    ROW0_DELAY    : in     std_logic_vector (abits_g-1 downto 0);
    PAGE_START    : in     std_logic_vector (25 downto 0);
    SYNC          : in     std_logic;
    CONV_ENABLE   : in     std_logic
  );

-- Declarations

end entity fop_str ;

