-- PCIE_HIP_FDAS.vhd

-- Generated using ACDS version 22.4 94

library IEEE;
library PCIE_HIP_FDAS_clock_bridge_0;
library PCIE_HIP_FDAS_mm_wr_transparent_0;
library PCIE_HIP_FDAS_mm_wr_transparent_1;
library PCIE_HIP_FDAS_mm_wr_transparent_2;
library PCIE_HIP_FDAS_mm_wr_transparent_3;
library PCIE_HIP_FDAS_mm_rd_transparent_0;
library PCIE_HIP_FDAS_mm_rd_transparent_1;
library PCIE_HIP_FDAS_mm_rd_transparent_2;
library PCIE_HIP_FDAS_mm_rd_transparent_3;
library PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0;
library PCIE_HIP_FDAS_reset_bridge_0;
library PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0;
library altera_mm_interconnect_1920;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PCIE_HIP_FDAS is
	port (
		clk_out_clk                                    : out std_logic;                                         --                              clk_out.clk
		rd_dma_0_waitrequest                           : in  std_logic                      := '0';             --                             rd_dma_0.waitrequest
		rd_dma_0_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		rd_dma_0_writedata                             : out std_logic_vector(511 downto 0);                    --                                     .writedata
		rd_dma_0_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		rd_dma_0_write                                 : out std_logic;                                         --                                     .write
		rd_dma_0_byteenable                            : out std_logic_vector(63 downto 0);                     --                                     .byteenable
		rd_dma_1_waitrequest                           : in  std_logic                      := '0';             --                             rd_dma_1.waitrequest
		rd_dma_1_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		rd_dma_1_writedata                             : out std_logic_vector(511 downto 0);                    --                                     .writedata
		rd_dma_1_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		rd_dma_1_write                                 : out std_logic;                                         --                                     .write
		rd_dma_1_byteenable                            : out std_logic_vector(63 downto 0);                     --                                     .byteenable
		rd_dma_2_waitrequest                           : in  std_logic                      := '0';             --                             rd_dma_2.waitrequest
		rd_dma_2_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		rd_dma_2_writedata                             : out std_logic_vector(511 downto 0);                    --                                     .writedata
		rd_dma_2_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		rd_dma_2_write                                 : out std_logic;                                         --                                     .write
		rd_dma_2_byteenable                            : out std_logic_vector(63 downto 0);                     --                                     .byteenable
		rd_dma_3_waitrequest                           : in  std_logic                      := '0';             --                             rd_dma_3.waitrequest
		rd_dma_3_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		rd_dma_3_writedata                             : out std_logic_vector(511 downto 0);                    --                                     .writedata
		rd_dma_3_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		rd_dma_3_write                                 : out std_logic;                                         --                                     .write
		rd_dma_3_byteenable                            : out std_logic_vector(63 downto 0);                     --                                     .byteenable
		wr_dma_0_waitrequest                           : in  std_logic                      := '0';             --                             wr_dma_0.waitrequest
		wr_dma_0_readdata                              : in  std_logic_vector(511 downto 0) := (others => '0'); --                                     .readdata
		wr_dma_0_readdatavalid                         : in  std_logic                      := '0';             --                                     .readdatavalid
		wr_dma_0_response                              : in  std_logic_vector(1 downto 0)   := (others => '0'); --                                     .response
		wr_dma_0_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		wr_dma_0_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		wr_dma_0_read                                  : out std_logic;                                         --                                     .read
		wr_dma_1_waitrequest                           : in  std_logic                      := '0';             --                             wr_dma_1.waitrequest
		wr_dma_1_readdata                              : in  std_logic_vector(511 downto 0) := (others => '0'); --                                     .readdata
		wr_dma_1_readdatavalid                         : in  std_logic                      := '0';             --                                     .readdatavalid
		wr_dma_1_response                              : in  std_logic_vector(1 downto 0)   := (others => '0'); --                                     .response
		wr_dma_1_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		wr_dma_1_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		wr_dma_1_read                                  : out std_logic;                                         --                                     .read
		wr_dma_2_waitrequest                           : in  std_logic                      := '0';             --                             wr_dma_2.waitrequest
		wr_dma_2_readdata                              : in  std_logic_vector(511 downto 0) := (others => '0'); --                                     .readdata
		wr_dma_2_readdatavalid                         : in  std_logic                      := '0';             --                                     .readdatavalid
		wr_dma_2_response                              : in  std_logic_vector(1 downto 0)   := (others => '0'); --                                     .response
		wr_dma_2_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		wr_dma_2_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		wr_dma_2_read                                  : out std_logic;                                         --                                     .read
		wr_dma_3_waitrequest                           : in  std_logic                      := '0';             --                             wr_dma_3.waitrequest
		wr_dma_3_readdata                              : in  std_logic_vector(511 downto 0) := (others => '0'); --                                     .readdata
		wr_dma_3_readdatavalid                         : in  std_logic                      := '0';             --                                     .readdatavalid
		wr_dma_3_response                              : in  std_logic_vector(1 downto 0)   := (others => '0'); --                                     .response
		wr_dma_3_burstcount                            : out std_logic_vector(3 downto 0);                      --                                     .burstcount
		wr_dma_3_address                               : out std_logic_vector(25 downto 0);                     --                                     .address
		wr_dma_3_read                                  : out std_logic;                                         --                                     .read
		intel_pcie_ptile_mcdma_0_p0_usr_msix_valid     : in  std_logic                      := '0';             -- intel_pcie_ptile_mcdma_0_p0_usr_msix.valid
		intel_pcie_ptile_mcdma_0_p0_usr_msix_ready     : out std_logic;                                         --                                     .ready
		intel_pcie_ptile_mcdma_0_p0_usr_msix_data      : in  std_logic_vector(15 downto 0)  := (others => '0'); --                                     .data
		intel_pcie_ptile_mcdma_0_refclk0_clk           : in  std_logic                      := '0';             --     intel_pcie_ptile_mcdma_0_refclk0.clk
		intel_pcie_ptile_mcdma_0_refclk1_clk           : in  std_logic                      := '0';             --     intel_pcie_ptile_mcdma_0_refclk1.clk
		intel_pcie_ptile_mcdma_0_ninit_done_reset      : in  std_logic                      := '0';             --  intel_pcie_ptile_mcdma_0_ninit_done.reset
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in0   : in  std_logic                      := '0';             --  intel_pcie_ptile_mcdma_0_hip_serial.rx_n_in0
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in1   : in  std_logic                      := '0';             --                                     .rx_n_in1
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in2   : in  std_logic                      := '0';             --                                     .rx_n_in2
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in3   : in  std_logic                      := '0';             --                                     .rx_n_in3
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in4   : in  std_logic                      := '0';             --                                     .rx_n_in4
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in5   : in  std_logic                      := '0';             --                                     .rx_n_in5
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in6   : in  std_logic                      := '0';             --                                     .rx_n_in6
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in7   : in  std_logic                      := '0';             --                                     .rx_n_in7
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in8   : in  std_logic                      := '0';             --                                     .rx_n_in8
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in9   : in  std_logic                      := '0';             --                                     .rx_n_in9
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in10  : in  std_logic                      := '0';             --                                     .rx_n_in10
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in11  : in  std_logic                      := '0';             --                                     .rx_n_in11
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in12  : in  std_logic                      := '0';             --                                     .rx_n_in12
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in13  : in  std_logic                      := '0';             --                                     .rx_n_in13
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in14  : in  std_logic                      := '0';             --                                     .rx_n_in14
		intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in15  : in  std_logic                      := '0';             --                                     .rx_n_in15
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in0   : in  std_logic                      := '0';             --                                     .rx_p_in0
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in1   : in  std_logic                      := '0';             --                                     .rx_p_in1
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in2   : in  std_logic                      := '0';             --                                     .rx_p_in2
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in3   : in  std_logic                      := '0';             --                                     .rx_p_in3
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in4   : in  std_logic                      := '0';             --                                     .rx_p_in4
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in5   : in  std_logic                      := '0';             --                                     .rx_p_in5
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in6   : in  std_logic                      := '0';             --                                     .rx_p_in6
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in7   : in  std_logic                      := '0';             --                                     .rx_p_in7
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in8   : in  std_logic                      := '0';             --                                     .rx_p_in8
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in9   : in  std_logic                      := '0';             --                                     .rx_p_in9
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in10  : in  std_logic                      := '0';             --                                     .rx_p_in10
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in11  : in  std_logic                      := '0';             --                                     .rx_p_in11
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in12  : in  std_logic                      := '0';             --                                     .rx_p_in12
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in13  : in  std_logic                      := '0';             --                                     .rx_p_in13
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in14  : in  std_logic                      := '0';             --                                     .rx_p_in14
		intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in15  : in  std_logic                      := '0';             --                                     .rx_p_in15
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out0  : out std_logic;                                         --                                     .tx_n_out0
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out1  : out std_logic;                                         --                                     .tx_n_out1
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out2  : out std_logic;                                         --                                     .tx_n_out2
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out3  : out std_logic;                                         --                                     .tx_n_out3
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out4  : out std_logic;                                         --                                     .tx_n_out4
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out5  : out std_logic;                                         --                                     .tx_n_out5
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out6  : out std_logic;                                         --                                     .tx_n_out6
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out7  : out std_logic;                                         --                                     .tx_n_out7
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out8  : out std_logic;                                         --                                     .tx_n_out8
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out9  : out std_logic;                                         --                                     .tx_n_out9
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out10 : out std_logic;                                         --                                     .tx_n_out10
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out11 : out std_logic;                                         --                                     .tx_n_out11
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out12 : out std_logic;                                         --                                     .tx_n_out12
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out13 : out std_logic;                                         --                                     .tx_n_out13
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out14 : out std_logic;                                         --                                     .tx_n_out14
		intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out15 : out std_logic;                                         --                                     .tx_n_out15
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out0  : out std_logic;                                         --                                     .tx_p_out0
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out1  : out std_logic;                                         --                                     .tx_p_out1
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out2  : out std_logic;                                         --                                     .tx_p_out2
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out3  : out std_logic;                                         --                                     .tx_p_out3
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out4  : out std_logic;                                         --                                     .tx_p_out4
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out5  : out std_logic;                                         --                                     .tx_p_out5
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out6  : out std_logic;                                         --                                     .tx_p_out6
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out7  : out std_logic;                                         --                                     .tx_p_out7
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out8  : out std_logic;                                         --                                     .tx_p_out8
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out9  : out std_logic;                                         --                                     .tx_p_out9
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out10 : out std_logic;                                         --                                     .tx_p_out10
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out11 : out std_logic;                                         --                                     .tx_p_out11
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out12 : out std_logic;                                         --                                     .tx_p_out12
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out13 : out std_logic;                                         --                                     .tx_p_out13
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out14 : out std_logic;                                         --                                     .tx_p_out14
		intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out15 : out std_logic;                                         --                                     .tx_p_out15
		intel_pcie_ptile_mcdma_0_pin_perst_reset_n     : in  std_logic                      := '0';             --   intel_pcie_ptile_mcdma_0_pin_perst.reset_n
		reset_out_reset_n                              : out std_logic;                                         --                            reset_out.reset_n
		rxm_bar2_0_m0_waitrequest                      : in  std_logic                      := '0';             --                        rxm_bar2_0_m0.waitrequest
		rxm_bar2_0_m0_readdata                         : in  std_logic_vector(63 downto 0)  := (others => '0'); --                                     .readdata
		rxm_bar2_0_m0_readdatavalid                    : in  std_logic                      := '0';             --                                     .readdatavalid
		rxm_bar2_0_m0_writeresponsevalid               : in  std_logic                      := '0';             --                                     .writeresponsevalid
		rxm_bar2_0_m0_response                         : in  std_logic_vector(1 downto 0)   := (others => '0'); --                                     .response
		rxm_bar2_0_m0_writedata                        : out std_logic_vector(63 downto 0);                     --                                     .writedata
		rxm_bar2_0_m0_address                          : out std_logic_vector(21 downto 0);                     --                                     .address
		rxm_bar2_0_m0_write                            : out std_logic;                                         --                                     .write
		rxm_bar2_0_m0_read                             : out std_logic;                                         --                                     .read
		rxm_bar2_0_m0_byteenable                       : out std_logic_vector(7 downto 0)                       --                                     .byteenable
	);
end entity PCIE_HIP_FDAS;

architecture rtl of PCIE_HIP_FDAS is
	component PCIE_HIP_FDAS_clock_bridge_0_cmp is
		port (
			in_clk  : in  std_logic := 'X'; -- clk
			out_clk : out std_logic         -- clk
		);
	end component PCIE_HIP_FDAS_clock_bridge_0_cmp;

	component PCIE_HIP_FDAS_mm_wr_transparent_0_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk            : in  std_logic                      := 'X';             -- clk
			reset          : in  std_logic                      := 'X';             -- reset
			s0_waitrequest : out std_logic;                                         -- waitrequest
			s0_burstcount  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_writedata   : in  std_logic_vector(511 downto 0) := (others => 'X'); -- writedata
			s0_address     : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_write       : in  std_logic                      := 'X';             -- write
			s0_byteenable  : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- byteenable
			m0_waitrequest : in  std_logic                      := 'X';             -- waitrequest
			m0_burstcount  : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_writedata   : out std_logic_vector(511 downto 0);                    -- writedata
			m0_address     : out std_logic_vector(25 downto 0);                     -- address
			m0_write       : out std_logic;                                         -- write
			m0_byteenable  : out std_logic_vector(63 downto 0)                      -- byteenable
		);
	end component PCIE_HIP_FDAS_mm_wr_transparent_0_cmp;

	component PCIE_HIP_FDAS_mm_wr_transparent_1_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk            : in  std_logic                      := 'X';             -- clk
			reset          : in  std_logic                      := 'X';             -- reset
			s0_waitrequest : out std_logic;                                         -- waitrequest
			s0_burstcount  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_writedata   : in  std_logic_vector(511 downto 0) := (others => 'X'); -- writedata
			s0_address     : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_write       : in  std_logic                      := 'X';             -- write
			s0_byteenable  : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- byteenable
			m0_waitrequest : in  std_logic                      := 'X';             -- waitrequest
			m0_burstcount  : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_writedata   : out std_logic_vector(511 downto 0);                    -- writedata
			m0_address     : out std_logic_vector(25 downto 0);                     -- address
			m0_write       : out std_logic;                                         -- write
			m0_byteenable  : out std_logic_vector(63 downto 0)                      -- byteenable
		);
	end component PCIE_HIP_FDAS_mm_wr_transparent_1_cmp;

	component PCIE_HIP_FDAS_mm_wr_transparent_2_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk            : in  std_logic                      := 'X';             -- clk
			reset          : in  std_logic                      := 'X';             -- reset
			s0_waitrequest : out std_logic;                                         -- waitrequest
			s0_burstcount  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_writedata   : in  std_logic_vector(511 downto 0) := (others => 'X'); -- writedata
			s0_address     : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_write       : in  std_logic                      := 'X';             -- write
			s0_byteenable  : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- byteenable
			m0_waitrequest : in  std_logic                      := 'X';             -- waitrequest
			m0_burstcount  : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_writedata   : out std_logic_vector(511 downto 0);                    -- writedata
			m0_address     : out std_logic_vector(25 downto 0);                     -- address
			m0_write       : out std_logic;                                         -- write
			m0_byteenable  : out std_logic_vector(63 downto 0)                      -- byteenable
		);
	end component PCIE_HIP_FDAS_mm_wr_transparent_2_cmp;

	component PCIE_HIP_FDAS_mm_wr_transparent_3_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk            : in  std_logic                      := 'X';             -- clk
			reset          : in  std_logic                      := 'X';             -- reset
			s0_waitrequest : out std_logic;                                         -- waitrequest
			s0_burstcount  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_writedata   : in  std_logic_vector(511 downto 0) := (others => 'X'); -- writedata
			s0_address     : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_write       : in  std_logic                      := 'X';             -- write
			s0_byteenable  : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- byteenable
			m0_waitrequest : in  std_logic                      := 'X';             -- waitrequest
			m0_burstcount  : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_writedata   : out std_logic_vector(511 downto 0);                    -- writedata
			m0_address     : out std_logic_vector(25 downto 0);                     -- address
			m0_write       : out std_logic;                                         -- write
			m0_byteenable  : out std_logic_vector(63 downto 0)                      -- byteenable
		);
	end component PCIE_HIP_FDAS_mm_wr_transparent_3_cmp;

	component PCIE_HIP_FDAS_mm_rd_transparent_0_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                         -- waitrequest
			s0_readdata      : out std_logic_vector(511 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                         -- readdatavalid
			s0_response      : out std_logic_vector(1 downto 0);                      -- response
			s0_burstcount    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_address       : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_read          : in  std_logic                      := 'X';             -- read
			m0_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			m0_response      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_burstcount    : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_address       : out std_logic_vector(25 downto 0);                     -- address
			m0_read          : out std_logic                                          -- read
		);
	end component PCIE_HIP_FDAS_mm_rd_transparent_0_cmp;

	component PCIE_HIP_FDAS_mm_rd_transparent_1_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                         -- waitrequest
			s0_readdata      : out std_logic_vector(511 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                         -- readdatavalid
			s0_response      : out std_logic_vector(1 downto 0);                      -- response
			s0_burstcount    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_address       : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_read          : in  std_logic                      := 'X';             -- read
			m0_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			m0_response      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_burstcount    : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_address       : out std_logic_vector(25 downto 0);                     -- address
			m0_read          : out std_logic                                          -- read
		);
	end component PCIE_HIP_FDAS_mm_rd_transparent_1_cmp;

	component PCIE_HIP_FDAS_mm_rd_transparent_2_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                         -- waitrequest
			s0_readdata      : out std_logic_vector(511 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                         -- readdatavalid
			s0_response      : out std_logic_vector(1 downto 0);                      -- response
			s0_burstcount    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_address       : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_read          : in  std_logic                      := 'X';             -- read
			m0_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			m0_response      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_burstcount    : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_address       : out std_logic_vector(25 downto 0);                     -- address
			m0_read          : out std_logic                                          -- read
		);
	end component PCIE_HIP_FDAS_mm_rd_transparent_2_cmp;

	component PCIE_HIP_FDAS_mm_rd_transparent_3_cmp is
		generic (
			DATA_WIDTH       : integer := 512;
			BYTE_SIZE        : integer := 8;
			ADDRESS_WIDTH    : integer := 26;
			BURSTCOUNT_WIDTH : integer := 4
		);
		port (
			clk              : in  std_logic                      := 'X';             -- clk
			reset            : in  std_logic                      := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                         -- waitrequest
			s0_readdata      : out std_logic_vector(511 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                         -- readdatavalid
			s0_response      : out std_logic_vector(1 downto 0);                      -- response
			s0_burstcount    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			s0_address       : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			s0_read          : in  std_logic                      := 'X';             -- read
			m0_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			m0_response      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_burstcount    : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_address       : out std_logic_vector(25 downto 0);                     -- address
			m0_read          : out std_logic                                          -- read
		);
	end component PCIE_HIP_FDAS_mm_rd_transparent_3_cmp;

	component PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0_cmp is
		port (
			app_clk                     : out std_logic;                                         -- clk
			app_rst_n                   : out std_logic;                                         -- reset_n
			rx_pio_waitrequest_i        : in  std_logic                      := 'X';             -- waitrequest
			rx_pio_address_o            : out std_logic_vector(27 downto 0);                     -- address
			rx_pio_byteenable_o         : out std_logic_vector(7 downto 0);                      -- byteenable
			rx_pio_read_o               : out std_logic;                                         -- read
			rx_pio_readdata_i           : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- readdata
			rx_pio_readdatavalid_i      : in  std_logic                      := 'X';             -- readdatavalid
			rx_pio_write_o              : out std_logic;                                         -- write
			rx_pio_writedata_o          : out std_logic_vector(63 downto 0);                     -- writedata
			rx_pio_burstcount_o         : out std_logic_vector(3 downto 0);                      -- burstcount
			rx_pio_response_i           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			rx_pio_writeresponsevalid_i : in  std_logic                      := 'X';             -- writeresponsevalid
			d2hdm_waitrequest_i         : in  std_logic                      := 'X';             -- waitrequest
			d2hdm_read_o                : out std_logic;                                         -- read
			d2hdm_address_o             : out std_logic_vector(63 downto 0);                     -- address
			d2hdm_burstcount_o          : out std_logic_vector(3 downto 0);                      -- burstcount
			d2hdm_byteenable_o          : out std_logic_vector(63 downto 0);                     -- byteenable
			d2hdm_readdatavalid_i       : in  std_logic                      := 'X';             -- readdatavalid
			d2hdm_readdata_i            : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			d2hdm_response_i            : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			h2ddm_waitrequest_i         : in  std_logic                      := 'X';             -- waitrequest
			h2ddm_write_o               : out std_logic;                                         -- write
			h2ddm_address_o             : out std_logic_vector(63 downto 0);                     -- address
			h2ddm_burstcount_o          : out std_logic_vector(3 downto 0);                      -- burstcount
			h2ddm_byteenable_o          : out std_logic_vector(63 downto 0);                     -- byteenable
			h2ddm_writedata_o           : out std_logic_vector(511 downto 0);                    -- writedata
			usr_event_msix_valid_i      : in  std_logic                      := 'X';             -- valid
			usr_event_msix_ready_o      : out std_logic;                                         -- ready
			usr_event_msix_data_i       : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- data
			usr_hip_tl_cfg_func_o       : out std_logic_vector(2 downto 0);                      -- tl_cfg_func
			usr_hip_tl_cfg_add_o        : out std_logic_vector(4 downto 0);                      -- tl_cfg_add
			usr_hip_tl_cfg_ctl_o        : out std_logic_vector(15 downto 0);                     -- tl_cfg_ctl
			p0_link_up_o                : out std_logic;                                         -- link_up
			p0_dl_up_o                  : out std_logic;                                         -- dl_up
			p0_surprise_down_err_o      : out std_logic;                                         -- surprise_down_err
			p0_ltssm_state_o            : out std_logic_vector(5 downto 0);                      -- ltssmstate
			refclk0                     : in  std_logic                      := 'X';             -- clk
			refclk1                     : in  std_logic                      := 'X';             -- clk
			ninit_done                  : in  std_logic                      := 'X';             -- reset
			rx_n_in0                    : in  std_logic                      := 'X';             -- rx_n_in0
			rx_n_in1                    : in  std_logic                      := 'X';             -- rx_n_in1
			rx_n_in2                    : in  std_logic                      := 'X';             -- rx_n_in2
			rx_n_in3                    : in  std_logic                      := 'X';             -- rx_n_in3
			rx_n_in4                    : in  std_logic                      := 'X';             -- rx_n_in4
			rx_n_in5                    : in  std_logic                      := 'X';             -- rx_n_in5
			rx_n_in6                    : in  std_logic                      := 'X';             -- rx_n_in6
			rx_n_in7                    : in  std_logic                      := 'X';             -- rx_n_in7
			rx_n_in8                    : in  std_logic                      := 'X';             -- rx_n_in8
			rx_n_in9                    : in  std_logic                      := 'X';             -- rx_n_in9
			rx_n_in10                   : in  std_logic                      := 'X';             -- rx_n_in10
			rx_n_in11                   : in  std_logic                      := 'X';             -- rx_n_in11
			rx_n_in12                   : in  std_logic                      := 'X';             -- rx_n_in12
			rx_n_in13                   : in  std_logic                      := 'X';             -- rx_n_in13
			rx_n_in14                   : in  std_logic                      := 'X';             -- rx_n_in14
			rx_n_in15                   : in  std_logic                      := 'X';             -- rx_n_in15
			rx_p_in0                    : in  std_logic                      := 'X';             -- rx_p_in0
			rx_p_in1                    : in  std_logic                      := 'X';             -- rx_p_in1
			rx_p_in2                    : in  std_logic                      := 'X';             -- rx_p_in2
			rx_p_in3                    : in  std_logic                      := 'X';             -- rx_p_in3
			rx_p_in4                    : in  std_logic                      := 'X';             -- rx_p_in4
			rx_p_in5                    : in  std_logic                      := 'X';             -- rx_p_in5
			rx_p_in6                    : in  std_logic                      := 'X';             -- rx_p_in6
			rx_p_in7                    : in  std_logic                      := 'X';             -- rx_p_in7
			rx_p_in8                    : in  std_logic                      := 'X';             -- rx_p_in8
			rx_p_in9                    : in  std_logic                      := 'X';             -- rx_p_in9
			rx_p_in10                   : in  std_logic                      := 'X';             -- rx_p_in10
			rx_p_in11                   : in  std_logic                      := 'X';             -- rx_p_in11
			rx_p_in12                   : in  std_logic                      := 'X';             -- rx_p_in12
			rx_p_in13                   : in  std_logic                      := 'X';             -- rx_p_in13
			rx_p_in14                   : in  std_logic                      := 'X';             -- rx_p_in14
			rx_p_in15                   : in  std_logic                      := 'X';             -- rx_p_in15
			tx_n_out0                   : out std_logic;                                         -- tx_n_out0
			tx_n_out1                   : out std_logic;                                         -- tx_n_out1
			tx_n_out2                   : out std_logic;                                         -- tx_n_out2
			tx_n_out3                   : out std_logic;                                         -- tx_n_out3
			tx_n_out4                   : out std_logic;                                         -- tx_n_out4
			tx_n_out5                   : out std_logic;                                         -- tx_n_out5
			tx_n_out6                   : out std_logic;                                         -- tx_n_out6
			tx_n_out7                   : out std_logic;                                         -- tx_n_out7
			tx_n_out8                   : out std_logic;                                         -- tx_n_out8
			tx_n_out9                   : out std_logic;                                         -- tx_n_out9
			tx_n_out10                  : out std_logic;                                         -- tx_n_out10
			tx_n_out11                  : out std_logic;                                         -- tx_n_out11
			tx_n_out12                  : out std_logic;                                         -- tx_n_out12
			tx_n_out13                  : out std_logic;                                         -- tx_n_out13
			tx_n_out14                  : out std_logic;                                         -- tx_n_out14
			tx_n_out15                  : out std_logic;                                         -- tx_n_out15
			tx_p_out0                   : out std_logic;                                         -- tx_p_out0
			tx_p_out1                   : out std_logic;                                         -- tx_p_out1
			tx_p_out2                   : out std_logic;                                         -- tx_p_out2
			tx_p_out3                   : out std_logic;                                         -- tx_p_out3
			tx_p_out4                   : out std_logic;                                         -- tx_p_out4
			tx_p_out5                   : out std_logic;                                         -- tx_p_out5
			tx_p_out6                   : out std_logic;                                         -- tx_p_out6
			tx_p_out7                   : out std_logic;                                         -- tx_p_out7
			tx_p_out8                   : out std_logic;                                         -- tx_p_out8
			tx_p_out9                   : out std_logic;                                         -- tx_p_out9
			tx_p_out10                  : out std_logic;                                         -- tx_p_out10
			tx_p_out11                  : out std_logic;                                         -- tx_p_out11
			tx_p_out12                  : out std_logic;                                         -- tx_p_out12
			tx_p_out13                  : out std_logic;                                         -- tx_p_out13
			tx_p_out14                  : out std_logic;                                         -- tx_p_out14
			tx_p_out15                  : out std_logic;                                         -- tx_p_out15
			pin_perst_n                 : in  std_logic                      := 'X'              -- reset_n
		);
	end component PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0_cmp;

	component PCIE_HIP_FDAS_reset_bridge_0_cmp is
		port (
			clk         : in  std_logic := 'X'; -- clk
			in_reset_n  : in  std_logic := 'X'; -- reset_n
			out_reset_n : out std_logic         -- reset_n
		);
	end component PCIE_HIP_FDAS_reset_bridge_0_cmp;

	component PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0_cmp is
		generic (
			DATA_WIDTH     : integer := 64;
			BYTE_SIZE      : integer := 8;
			ADDRESS_WIDTH  : integer := 22;
			RESPONSE_WIDTH : integer := 2
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			s0_waitrequest        : out std_logic;                                        -- waitrequest
			s0_readdata           : out std_logic_vector(63 downto 0);                    -- readdata
			s0_readdatavalid      : out std_logic;                                        -- readdatavalid
			s0_writeresponsevalid : out std_logic;                                        -- writeresponsevalid
			s0_response           : out std_logic_vector(1 downto 0);                     -- response
			s0_writedata          : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			s0_address            : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			s0_write              : in  std_logic                     := 'X';             -- write
			s0_read               : in  std_logic                     := 'X';             -- read
			s0_byteenable         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			m0_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata           : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			m0_writeresponsevalid : in  std_logic                     := 'X';             -- writeresponsevalid
			m0_response           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writedata          : out std_logic_vector(63 downto 0);                    -- writedata
			m0_address            : out std_logic_vector(21 downto 0);                    -- address
			m0_write              : out std_logic;                                        -- write
			m0_read               : out std_logic;                                        -- read
			m0_byteenable         : out std_logic_vector(7 downto 0)                      -- byteenable
		);
	end component PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0_cmp;

	component PCIE_HIP_FDAS_altera_mm_interconnect_1920_yasd64i_cmp is
		port (
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_address                                      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_waitrequest                                  : out std_logic;                                         -- waitrequest
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_burstcount                                   : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_byteenable                                   : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- byteenable
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_read                                         : in  std_logic                      := 'X';             -- read
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdata                                     : out std_logic_vector(511 downto 0);                    -- readdata
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdatavalid                                : out std_logic;                                         -- readdatavalid
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_response                                     : out std_logic_vector(1 downto 0);                      -- response
			dma_wr_0_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_wr_0_s0_read                                                                      : out std_logic;                                         -- read
			dma_wr_0_s0_readdata                                                                  : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			dma_wr_0_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_wr_0_s0_readdatavalid                                                             : in  std_logic                      := 'X';             -- readdatavalid
			dma_wr_0_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_wr_0_s0_response                                                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			dma_wr_1_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_wr_1_s0_read                                                                      : out std_logic;                                         -- read
			dma_wr_1_s0_readdata                                                                  : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			dma_wr_1_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_wr_1_s0_readdatavalid                                                             : in  std_logic                      := 'X';             -- readdatavalid
			dma_wr_1_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_wr_1_s0_response                                                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			dma_wr_2_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_wr_2_s0_read                                                                      : out std_logic;                                         -- read
			dma_wr_2_s0_readdata                                                                  : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			dma_wr_2_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_wr_2_s0_readdatavalid                                                             : in  std_logic                      := 'X';             -- readdatavalid
			dma_wr_2_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_wr_2_s0_response                                                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			dma_wr_3_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_wr_3_s0_read                                                                      : out std_logic;                                         -- read
			dma_wr_3_s0_readdata                                                                  : in  std_logic_vector(511 downto 0) := (others => 'X'); -- readdata
			dma_wr_3_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_wr_3_s0_readdatavalid                                                             : in  std_logic                      := 'X';             -- readdatavalid
			dma_wr_3_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_wr_3_s0_response                                                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			dma_wr_0_reset_reset_bridge_in_reset_reset                                            : in  std_logic                      := 'X';             -- reset
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			intel_pcie_ptile_mcdma_0_app_clk_clk                                                  : in  std_logic                      := 'X'              -- clk
		);
	end component PCIE_HIP_FDAS_altera_mm_interconnect_1920_yasd64i_cmp;

	component PCIE_HIP_FDAS_altera_mm_interconnect_1920_j3desai_cmp is
		port (
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_address                                      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_waitrequest                                  : out std_logic;                                         -- waitrequest
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_burstcount                                   : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_byteenable                                   : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- byteenable
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_write                                        : in  std_logic                      := 'X';             -- write
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_writedata                                    : in  std_logic_vector(511 downto 0) := (others => 'X'); -- writedata
			dma_rd_0_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_rd_0_s0_write                                                                     : out std_logic;                                         -- write
			dma_rd_0_s0_writedata                                                                 : out std_logic_vector(511 downto 0);                    -- writedata
			dma_rd_0_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_rd_0_s0_byteenable                                                                : out std_logic_vector(63 downto 0);                     -- byteenable
			dma_rd_0_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_rd_1_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_rd_1_s0_write                                                                     : out std_logic;                                         -- write
			dma_rd_1_s0_writedata                                                                 : out std_logic_vector(511 downto 0);                    -- writedata
			dma_rd_1_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_rd_1_s0_byteenable                                                                : out std_logic_vector(63 downto 0);                     -- byteenable
			dma_rd_1_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_rd_2_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_rd_2_s0_write                                                                     : out std_logic;                                         -- write
			dma_rd_2_s0_writedata                                                                 : out std_logic_vector(511 downto 0);                    -- writedata
			dma_rd_2_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_rd_2_s0_byteenable                                                                : out std_logic_vector(63 downto 0);                     -- byteenable
			dma_rd_2_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_rd_3_s0_address                                                                   : out std_logic_vector(25 downto 0);                     -- address
			dma_rd_3_s0_write                                                                     : out std_logic;                                         -- write
			dma_rd_3_s0_writedata                                                                 : out std_logic_vector(511 downto 0);                    -- writedata
			dma_rd_3_s0_burstcount                                                                : out std_logic_vector(3 downto 0);                      -- burstcount
			dma_rd_3_s0_byteenable                                                                : out std_logic_vector(63 downto 0);                     -- byteenable
			dma_rd_3_s0_waitrequest                                                               : in  std_logic                      := 'X';             -- waitrequest
			dma_rd_0_reset_reset_bridge_in_reset_reset                                            : in  std_logic                      := 'X';             -- reset
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			intel_pcie_ptile_mcdma_0_app_clk_clk                                                  : in  std_logic                      := 'X'              -- clk
		);
	end component PCIE_HIP_FDAS_altera_mm_interconnect_1920_j3desai_cmp;

	component PCIE_HIP_FDAS_altera_mm_interconnect_1920_jrv6pua_cmp is
		port (
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_address                                      : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_waitrequest                                  : out std_logic;                                        -- waitrequest
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_burstcount                                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_byteenable                                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_read                                         : in  std_logic                     := 'X';             -- read
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdata                                     : out std_logic_vector(63 downto 0);                    -- readdata
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdatavalid                                : out std_logic;                                        -- readdatavalid
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_write                                        : in  std_logic                     := 'X';             -- write
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writedata                                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_response                                     : out std_logic_vector(1 downto 0);                     -- response
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writeresponsevalid                           : out std_logic;                                        -- writeresponsevalid
			rxm_bar2_0_s0_address                                                                  : out std_logic_vector(21 downto 0);                    -- address
			rxm_bar2_0_s0_write                                                                    : out std_logic;                                        -- write
			rxm_bar2_0_s0_read                                                                     : out std_logic;                                        -- read
			rxm_bar2_0_s0_readdata                                                                 : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			rxm_bar2_0_s0_writedata                                                                : out std_logic_vector(63 downto 0);                    -- writedata
			rxm_bar2_0_s0_byteenable                                                               : out std_logic_vector(7 downto 0);                     -- byteenable
			rxm_bar2_0_s0_readdatavalid                                                            : in  std_logic                     := 'X';             -- readdatavalid
			rxm_bar2_0_s0_waitrequest                                                              : in  std_logic                     := 'X';             -- waitrequest
			rxm_bar2_0_s0_response                                                                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			rxm_bar2_0_s0_writeresponsevalid                                                       : in  std_logic                     := 'X';             -- writeresponsevalid
			rxm_bar2_0_reset_reset_bridge_in_reset_reset                                           : in  std_logic                     := 'X';             -- reset
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			intel_pcie_ptile_mcdma_0_app_clk_clk                                                   : in  std_logic                     := 'X'              -- clk
		);
	end component PCIE_HIP_FDAS_altera_mm_interconnect_1920_jrv6pua_cmp;

	signal intel_pcie_ptile_mcdma_0_app_clk_clk                         : std_logic;                      -- intel_pcie_ptile_mcdma_0:app_clk -> [clock_bridge_0:in_clk, dma_rd_0:clk, dma_rd_1:clk, dma_rd_2:clk, dma_rd_3:clk, dma_wr_0:clk, dma_wr_1:clk, dma_wr_2:clk, dma_wr_3:clk, mm_interconnect_0:intel_pcie_ptile_mcdma_0_app_clk_clk, mm_interconnect_1:intel_pcie_ptile_mcdma_0_app_clk_clk, mm_interconnect_2:intel_pcie_ptile_mcdma_0_app_clk_clk, reset_bridge_0:clk, rxm_bar2_0:clk]
	signal intel_pcie_ptile_mcdma_0_app_nreset_status_reset             : std_logic;                      -- intel_pcie_ptile_mcdma_0:app_rst_n -> [intel_pcie_ptile_mcdma_0_app_nreset_status_reset:in, reset_bridge_0:in_reset_n]
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_waitrequest         : std_logic;                      -- mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_waitrequest -> intel_pcie_ptile_mcdma_0:d2hdm_waitrequest_i
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdata            : std_logic_vector(511 downto 0); -- mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdata -> intel_pcie_ptile_mcdma_0:d2hdm_readdata_i
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_read                : std_logic;                      -- intel_pcie_ptile_mcdma_0:d2hdm_read_o -> mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_read
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_address             : std_logic_vector(63 downto 0);  -- intel_pcie_ptile_mcdma_0:d2hdm_address_o -> mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_address
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_byteenable          : std_logic_vector(63 downto 0);  -- intel_pcie_ptile_mcdma_0:d2hdm_byteenable_o -> mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_byteenable
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdatavalid       : std_logic;                      -- mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdatavalid -> intel_pcie_ptile_mcdma_0:d2hdm_readdatavalid_i
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_response            : std_logic_vector(1 downto 0);   -- mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_response -> intel_pcie_ptile_mcdma_0:d2hdm_response_i
	signal intel_pcie_ptile_mcdma_0_p0_d2hdm_master_burstcount          : std_logic_vector(3 downto 0);   -- intel_pcie_ptile_mcdma_0:d2hdm_burstcount_o -> mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_burstcount
	signal mm_interconnect_0_dma_wr_0_s0_readdata                       : std_logic_vector(511 downto 0); -- dma_wr_0:s0_readdata -> mm_interconnect_0:dma_wr_0_s0_readdata
	signal mm_interconnect_0_dma_wr_0_s0_waitrequest                    : std_logic;                      -- dma_wr_0:s0_waitrequest -> mm_interconnect_0:dma_wr_0_s0_waitrequest
	signal mm_interconnect_0_dma_wr_0_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_0:dma_wr_0_s0_address -> dma_wr_0:s0_address
	signal mm_interconnect_0_dma_wr_0_s0_read                           : std_logic;                      -- mm_interconnect_0:dma_wr_0_s0_read -> dma_wr_0:s0_read
	signal mm_interconnect_0_dma_wr_0_s0_readdatavalid                  : std_logic;                      -- dma_wr_0:s0_readdatavalid -> mm_interconnect_0:dma_wr_0_s0_readdatavalid
	signal mm_interconnect_0_dma_wr_0_s0_response                       : std_logic_vector(1 downto 0);   -- dma_wr_0:s0_response -> mm_interconnect_0:dma_wr_0_s0_response
	signal mm_interconnect_0_dma_wr_0_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_0:dma_wr_0_s0_burstcount -> dma_wr_0:s0_burstcount
	signal mm_interconnect_0_dma_wr_1_s0_readdata                       : std_logic_vector(511 downto 0); -- dma_wr_1:s0_readdata -> mm_interconnect_0:dma_wr_1_s0_readdata
	signal mm_interconnect_0_dma_wr_1_s0_waitrequest                    : std_logic;                      -- dma_wr_1:s0_waitrequest -> mm_interconnect_0:dma_wr_1_s0_waitrequest
	signal mm_interconnect_0_dma_wr_1_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_0:dma_wr_1_s0_address -> dma_wr_1:s0_address
	signal mm_interconnect_0_dma_wr_1_s0_read                           : std_logic;                      -- mm_interconnect_0:dma_wr_1_s0_read -> dma_wr_1:s0_read
	signal mm_interconnect_0_dma_wr_1_s0_readdatavalid                  : std_logic;                      -- dma_wr_1:s0_readdatavalid -> mm_interconnect_0:dma_wr_1_s0_readdatavalid
	signal mm_interconnect_0_dma_wr_1_s0_response                       : std_logic_vector(1 downto 0);   -- dma_wr_1:s0_response -> mm_interconnect_0:dma_wr_1_s0_response
	signal mm_interconnect_0_dma_wr_1_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_0:dma_wr_1_s0_burstcount -> dma_wr_1:s0_burstcount
	signal mm_interconnect_0_dma_wr_2_s0_readdata                       : std_logic_vector(511 downto 0); -- dma_wr_2:s0_readdata -> mm_interconnect_0:dma_wr_2_s0_readdata
	signal mm_interconnect_0_dma_wr_2_s0_waitrequest                    : std_logic;                      -- dma_wr_2:s0_waitrequest -> mm_interconnect_0:dma_wr_2_s0_waitrequest
	signal mm_interconnect_0_dma_wr_2_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_0:dma_wr_2_s0_address -> dma_wr_2:s0_address
	signal mm_interconnect_0_dma_wr_2_s0_read                           : std_logic;                      -- mm_interconnect_0:dma_wr_2_s0_read -> dma_wr_2:s0_read
	signal mm_interconnect_0_dma_wr_2_s0_readdatavalid                  : std_logic;                      -- dma_wr_2:s0_readdatavalid -> mm_interconnect_0:dma_wr_2_s0_readdatavalid
	signal mm_interconnect_0_dma_wr_2_s0_response                       : std_logic_vector(1 downto 0);   -- dma_wr_2:s0_response -> mm_interconnect_0:dma_wr_2_s0_response
	signal mm_interconnect_0_dma_wr_2_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_0:dma_wr_2_s0_burstcount -> dma_wr_2:s0_burstcount
	signal mm_interconnect_0_dma_wr_3_s0_readdata                       : std_logic_vector(511 downto 0); -- dma_wr_3:s0_readdata -> mm_interconnect_0:dma_wr_3_s0_readdata
	signal mm_interconnect_0_dma_wr_3_s0_waitrequest                    : std_logic;                      -- dma_wr_3:s0_waitrequest -> mm_interconnect_0:dma_wr_3_s0_waitrequest
	signal mm_interconnect_0_dma_wr_3_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_0:dma_wr_3_s0_address -> dma_wr_3:s0_address
	signal mm_interconnect_0_dma_wr_3_s0_read                           : std_logic;                      -- mm_interconnect_0:dma_wr_3_s0_read -> dma_wr_3:s0_read
	signal mm_interconnect_0_dma_wr_3_s0_readdatavalid                  : std_logic;                      -- dma_wr_3:s0_readdatavalid -> mm_interconnect_0:dma_wr_3_s0_readdatavalid
	signal mm_interconnect_0_dma_wr_3_s0_response                       : std_logic_vector(1 downto 0);   -- dma_wr_3:s0_response -> mm_interconnect_0:dma_wr_3_s0_response
	signal mm_interconnect_0_dma_wr_3_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_0:dma_wr_3_s0_burstcount -> dma_wr_3:s0_burstcount
	signal intel_pcie_ptile_mcdma_0_p0_h2ddm_master_waitrequest         : std_logic;                      -- mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_waitrequest -> intel_pcie_ptile_mcdma_0:h2ddm_waitrequest_i
	signal intel_pcie_ptile_mcdma_0_p0_h2ddm_master_address             : std_logic_vector(63 downto 0);  -- intel_pcie_ptile_mcdma_0:h2ddm_address_o -> mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_address
	signal intel_pcie_ptile_mcdma_0_p0_h2ddm_master_byteenable          : std_logic_vector(63 downto 0);  -- intel_pcie_ptile_mcdma_0:h2ddm_byteenable_o -> mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_byteenable
	signal intel_pcie_ptile_mcdma_0_p0_h2ddm_master_write               : std_logic;                      -- intel_pcie_ptile_mcdma_0:h2ddm_write_o -> mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_write
	signal intel_pcie_ptile_mcdma_0_p0_h2ddm_master_writedata           : std_logic_vector(511 downto 0); -- intel_pcie_ptile_mcdma_0:h2ddm_writedata_o -> mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_writedata
	signal intel_pcie_ptile_mcdma_0_p0_h2ddm_master_burstcount          : std_logic_vector(3 downto 0);   -- intel_pcie_ptile_mcdma_0:h2ddm_burstcount_o -> mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_burstcount
	signal mm_interconnect_1_dma_rd_0_s0_waitrequest                    : std_logic;                      -- dma_rd_0:s0_waitrequest -> mm_interconnect_1:dma_rd_0_s0_waitrequest
	signal mm_interconnect_1_dma_rd_0_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_1:dma_rd_0_s0_address -> dma_rd_0:s0_address
	signal mm_interconnect_1_dma_rd_0_s0_byteenable                     : std_logic_vector(63 downto 0);  -- mm_interconnect_1:dma_rd_0_s0_byteenable -> dma_rd_0:s0_byteenable
	signal mm_interconnect_1_dma_rd_0_s0_write                          : std_logic;                      -- mm_interconnect_1:dma_rd_0_s0_write -> dma_rd_0:s0_write
	signal mm_interconnect_1_dma_rd_0_s0_writedata                      : std_logic_vector(511 downto 0); -- mm_interconnect_1:dma_rd_0_s0_writedata -> dma_rd_0:s0_writedata
	signal mm_interconnect_1_dma_rd_0_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_rd_0_s0_burstcount -> dma_rd_0:s0_burstcount
	signal mm_interconnect_1_dma_rd_1_s0_waitrequest                    : std_logic;                      -- dma_rd_1:s0_waitrequest -> mm_interconnect_1:dma_rd_1_s0_waitrequest
	signal mm_interconnect_1_dma_rd_1_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_1:dma_rd_1_s0_address -> dma_rd_1:s0_address
	signal mm_interconnect_1_dma_rd_1_s0_byteenable                     : std_logic_vector(63 downto 0);  -- mm_interconnect_1:dma_rd_1_s0_byteenable -> dma_rd_1:s0_byteenable
	signal mm_interconnect_1_dma_rd_1_s0_write                          : std_logic;                      -- mm_interconnect_1:dma_rd_1_s0_write -> dma_rd_1:s0_write
	signal mm_interconnect_1_dma_rd_1_s0_writedata                      : std_logic_vector(511 downto 0); -- mm_interconnect_1:dma_rd_1_s0_writedata -> dma_rd_1:s0_writedata
	signal mm_interconnect_1_dma_rd_1_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_rd_1_s0_burstcount -> dma_rd_1:s0_burstcount
	signal mm_interconnect_1_dma_rd_2_s0_waitrequest                    : std_logic;                      -- dma_rd_2:s0_waitrequest -> mm_interconnect_1:dma_rd_2_s0_waitrequest
	signal mm_interconnect_1_dma_rd_2_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_1:dma_rd_2_s0_address -> dma_rd_2:s0_address
	signal mm_interconnect_1_dma_rd_2_s0_byteenable                     : std_logic_vector(63 downto 0);  -- mm_interconnect_1:dma_rd_2_s0_byteenable -> dma_rd_2:s0_byteenable
	signal mm_interconnect_1_dma_rd_2_s0_write                          : std_logic;                      -- mm_interconnect_1:dma_rd_2_s0_write -> dma_rd_2:s0_write
	signal mm_interconnect_1_dma_rd_2_s0_writedata                      : std_logic_vector(511 downto 0); -- mm_interconnect_1:dma_rd_2_s0_writedata -> dma_rd_2:s0_writedata
	signal mm_interconnect_1_dma_rd_2_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_rd_2_s0_burstcount -> dma_rd_2:s0_burstcount
	signal mm_interconnect_1_dma_rd_3_s0_waitrequest                    : std_logic;                      -- dma_rd_3:s0_waitrequest -> mm_interconnect_1:dma_rd_3_s0_waitrequest
	signal mm_interconnect_1_dma_rd_3_s0_address                        : std_logic_vector(25 downto 0);  -- mm_interconnect_1:dma_rd_3_s0_address -> dma_rd_3:s0_address
	signal mm_interconnect_1_dma_rd_3_s0_byteenable                     : std_logic_vector(63 downto 0);  -- mm_interconnect_1:dma_rd_3_s0_byteenable -> dma_rd_3:s0_byteenable
	signal mm_interconnect_1_dma_rd_3_s0_write                          : std_logic;                      -- mm_interconnect_1:dma_rd_3_s0_write -> dma_rd_3:s0_write
	signal mm_interconnect_1_dma_rd_3_s0_writedata                      : std_logic_vector(511 downto 0); -- mm_interconnect_1:dma_rd_3_s0_writedata -> dma_rd_3:s0_writedata
	signal mm_interconnect_1_dma_rd_3_s0_burstcount                     : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_rd_3_s0_burstcount -> dma_rd_3:s0_burstcount
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_waitrequest        : std_logic;                      -- mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_waitrequest -> intel_pcie_ptile_mcdma_0:rx_pio_waitrequest_i
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdata           : std_logic_vector(63 downto 0);  -- mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdata -> intel_pcie_ptile_mcdma_0:rx_pio_readdata_i
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_address            : std_logic_vector(27 downto 0);  -- intel_pcie_ptile_mcdma_0:rx_pio_address_o -> mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_address
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_byteenable         : std_logic_vector(7 downto 0);   -- intel_pcie_ptile_mcdma_0:rx_pio_byteenable_o -> mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_byteenable
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_read               : std_logic;                      -- intel_pcie_ptile_mcdma_0:rx_pio_read_o -> mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_read
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdatavalid      : std_logic;                      -- mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdatavalid -> intel_pcie_ptile_mcdma_0:rx_pio_readdatavalid_i
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_response           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_response -> intel_pcie_ptile_mcdma_0:rx_pio_response_i
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_write              : std_logic;                      -- intel_pcie_ptile_mcdma_0:rx_pio_write_o -> mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_write
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writedata          : std_logic_vector(63 downto 0);  -- intel_pcie_ptile_mcdma_0:rx_pio_writedata_o -> mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writedata
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writeresponsevalid : std_logic;                      -- mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writeresponsevalid -> intel_pcie_ptile_mcdma_0:rx_pio_writeresponsevalid_i
	signal intel_pcie_ptile_mcdma_0_p0_rx_pio_master_burstcount         : std_logic_vector(3 downto 0);   -- intel_pcie_ptile_mcdma_0:rx_pio_burstcount_o -> mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_burstcount
	signal mm_interconnect_2_rxm_bar2_0_s0_readdata                     : std_logic_vector(63 downto 0);  -- rxm_bar2_0:s0_readdata -> mm_interconnect_2:rxm_bar2_0_s0_readdata
	signal mm_interconnect_2_rxm_bar2_0_s0_waitrequest                  : std_logic;                      -- rxm_bar2_0:s0_waitrequest -> mm_interconnect_2:rxm_bar2_0_s0_waitrequest
	signal mm_interconnect_2_rxm_bar2_0_s0_address                      : std_logic_vector(21 downto 0);  -- mm_interconnect_2:rxm_bar2_0_s0_address -> rxm_bar2_0:s0_address
	signal mm_interconnect_2_rxm_bar2_0_s0_read                         : std_logic;                      -- mm_interconnect_2:rxm_bar2_0_s0_read -> rxm_bar2_0:s0_read
	signal mm_interconnect_2_rxm_bar2_0_s0_byteenable                   : std_logic_vector(7 downto 0);   -- mm_interconnect_2:rxm_bar2_0_s0_byteenable -> rxm_bar2_0:s0_byteenable
	signal mm_interconnect_2_rxm_bar2_0_s0_readdatavalid                : std_logic;                      -- rxm_bar2_0:s0_readdatavalid -> mm_interconnect_2:rxm_bar2_0_s0_readdatavalid
	signal mm_interconnect_2_rxm_bar2_0_s0_response                     : std_logic_vector(1 downto 0);   -- rxm_bar2_0:s0_response -> mm_interconnect_2:rxm_bar2_0_s0_response
	signal mm_interconnect_2_rxm_bar2_0_s0_write                        : std_logic;                      -- mm_interconnect_2:rxm_bar2_0_s0_write -> rxm_bar2_0:s0_write
	signal mm_interconnect_2_rxm_bar2_0_s0_writedata                    : std_logic_vector(63 downto 0);  -- mm_interconnect_2:rxm_bar2_0_s0_writedata -> rxm_bar2_0:s0_writedata
	signal mm_interconnect_2_rxm_bar2_0_s0_writeresponsevalid           : std_logic;                      -- rxm_bar2_0:s0_writeresponsevalid -> mm_interconnect_2:rxm_bar2_0_s0_writeresponsevalid
	signal intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv   : std_logic;                      -- intel_pcie_ptile_mcdma_0_app_nreset_status_reset:inv -> [dma_rd_0:reset, dma_rd_1:reset, dma_rd_2:reset, dma_rd_3:reset, dma_wr_0:reset, dma_wr_1:reset, dma_wr_2:reset, dma_wr_3:reset, mm_interconnect_0:dma_wr_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:intel_pcie_ptile_mcdma_0_p0_d2hdm_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:dma_rd_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:intel_pcie_ptile_mcdma_0_p0_h2ddm_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:intel_pcie_ptile_mcdma_0_p0_rx_pio_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:rxm_bar2_0_reset_reset_bridge_in_reset_reset, rxm_bar2_0:reset]

	for clock_bridge_0 : PCIE_HIP_FDAS_clock_bridge_0_cmp
		use entity PCIE_HIP_FDAS_clock_bridge_0.PCIE_HIP_FDAS_clock_bridge_0;
	for dma_rd_0 : PCIE_HIP_FDAS_mm_wr_transparent_0_cmp
		use entity PCIE_HIP_FDAS_mm_wr_transparent_0.PCIE_HIP_FDAS_mm_wr_transparent_0;
	for dma_rd_1 : PCIE_HIP_FDAS_mm_wr_transparent_1_cmp
		use entity PCIE_HIP_FDAS_mm_wr_transparent_1.PCIE_HIP_FDAS_mm_wr_transparent_1;
	for dma_rd_2 : PCIE_HIP_FDAS_mm_wr_transparent_2_cmp
		use entity PCIE_HIP_FDAS_mm_wr_transparent_2.PCIE_HIP_FDAS_mm_wr_transparent_2;
	for dma_rd_3 : PCIE_HIP_FDAS_mm_wr_transparent_3_cmp
		use entity PCIE_HIP_FDAS_mm_wr_transparent_3.PCIE_HIP_FDAS_mm_wr_transparent_3;
	for dma_wr_0 : PCIE_HIP_FDAS_mm_rd_transparent_0_cmp
		use entity PCIE_HIP_FDAS_mm_rd_transparent_0.PCIE_HIP_FDAS_mm_rd_transparent_0;
	for dma_wr_1 : PCIE_HIP_FDAS_mm_rd_transparent_1_cmp
		use entity PCIE_HIP_FDAS_mm_rd_transparent_1.PCIE_HIP_FDAS_mm_rd_transparent_1;
	for dma_wr_2 : PCIE_HIP_FDAS_mm_rd_transparent_2_cmp
		use entity PCIE_HIP_FDAS_mm_rd_transparent_2.PCIE_HIP_FDAS_mm_rd_transparent_2;
	for dma_wr_3 : PCIE_HIP_FDAS_mm_rd_transparent_3_cmp
		use entity PCIE_HIP_FDAS_mm_rd_transparent_3.PCIE_HIP_FDAS_mm_rd_transparent_3;
	for intel_pcie_ptile_mcdma_0 : PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0_cmp
		use entity PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0.PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0;
	for reset_bridge_0 : PCIE_HIP_FDAS_reset_bridge_0_cmp
		use entity PCIE_HIP_FDAS_reset_bridge_0.PCIE_HIP_FDAS_reset_bridge_0;
	for rxm_bar2_0 : PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0_cmp
		use entity PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0.PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0;
	for mm_interconnect_0 : PCIE_HIP_FDAS_altera_mm_interconnect_1920_yasd64i_cmp
		use entity altera_mm_interconnect_1920.PCIE_HIP_FDAS_altera_mm_interconnect_1920_yasd64i;
	for mm_interconnect_1 : PCIE_HIP_FDAS_altera_mm_interconnect_1920_j3desai_cmp
		use entity altera_mm_interconnect_1920.PCIE_HIP_FDAS_altera_mm_interconnect_1920_j3desai;
	for mm_interconnect_2 : PCIE_HIP_FDAS_altera_mm_interconnect_1920_jrv6pua_cmp
		use entity altera_mm_interconnect_1920.PCIE_HIP_FDAS_altera_mm_interconnect_1920_jrv6pua;
begin

	clock_bridge_0 : component PCIE_HIP_FDAS_clock_bridge_0_cmp
		port map (
			in_clk  => intel_pcie_ptile_mcdma_0_app_clk_clk, --  in_clk.clk
			out_clk => clk_out_clk                           -- out_clk.clk
		);

	dma_rd_0 : component PCIE_HIP_FDAS_mm_wr_transparent_0_cmp
		port map (
			clk            => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset          => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest => mm_interconnect_1_dma_rd_0_s0_waitrequest,                  --    s0.waitrequest
			s0_burstcount  => mm_interconnect_1_dma_rd_0_s0_burstcount,                   --      .burstcount
			s0_writedata   => mm_interconnect_1_dma_rd_0_s0_writedata,                    --      .writedata
			s0_address     => mm_interconnect_1_dma_rd_0_s0_address,                      --      .address
			s0_write       => mm_interconnect_1_dma_rd_0_s0_write,                        --      .write
			s0_byteenable  => mm_interconnect_1_dma_rd_0_s0_byteenable,                   --      .byteenable
			m0_waitrequest => rd_dma_0_waitrequest,                                       --    m0.waitrequest
			m0_burstcount  => rd_dma_0_burstcount,                                        --      .burstcount
			m0_writedata   => rd_dma_0_writedata,                                         --      .writedata
			m0_address     => rd_dma_0_address,                                           --      .address
			m0_write       => rd_dma_0_write,                                             --      .write
			m0_byteenable  => rd_dma_0_byteenable                                         --      .byteenable
		);

	dma_rd_1 : component PCIE_HIP_FDAS_mm_wr_transparent_1_cmp
		port map (
			clk            => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset          => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest => mm_interconnect_1_dma_rd_1_s0_waitrequest,                  --    s0.waitrequest
			s0_burstcount  => mm_interconnect_1_dma_rd_1_s0_burstcount,                   --      .burstcount
			s0_writedata   => mm_interconnect_1_dma_rd_1_s0_writedata,                    --      .writedata
			s0_address     => mm_interconnect_1_dma_rd_1_s0_address,                      --      .address
			s0_write       => mm_interconnect_1_dma_rd_1_s0_write,                        --      .write
			s0_byteenable  => mm_interconnect_1_dma_rd_1_s0_byteenable,                   --      .byteenable
			m0_waitrequest => rd_dma_1_waitrequest,                                       --    m0.waitrequest
			m0_burstcount  => rd_dma_1_burstcount,                                        --      .burstcount
			m0_writedata   => rd_dma_1_writedata,                                         --      .writedata
			m0_address     => rd_dma_1_address,                                           --      .address
			m0_write       => rd_dma_1_write,                                             --      .write
			m0_byteenable  => rd_dma_1_byteenable                                         --      .byteenable
		);

	dma_rd_2 : component PCIE_HIP_FDAS_mm_wr_transparent_2_cmp
		port map (
			clk            => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset          => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest => mm_interconnect_1_dma_rd_2_s0_waitrequest,                  --    s0.waitrequest
			s0_burstcount  => mm_interconnect_1_dma_rd_2_s0_burstcount,                   --      .burstcount
			s0_writedata   => mm_interconnect_1_dma_rd_2_s0_writedata,                    --      .writedata
			s0_address     => mm_interconnect_1_dma_rd_2_s0_address,                      --      .address
			s0_write       => mm_interconnect_1_dma_rd_2_s0_write,                        --      .write
			s0_byteenable  => mm_interconnect_1_dma_rd_2_s0_byteenable,                   --      .byteenable
			m0_waitrequest => rd_dma_2_waitrequest,                                       --    m0.waitrequest
			m0_burstcount  => rd_dma_2_burstcount,                                        --      .burstcount
			m0_writedata   => rd_dma_2_writedata,                                         --      .writedata
			m0_address     => rd_dma_2_address,                                           --      .address
			m0_write       => rd_dma_2_write,                                             --      .write
			m0_byteenable  => rd_dma_2_byteenable                                         --      .byteenable
		);

	dma_rd_3 : component PCIE_HIP_FDAS_mm_wr_transparent_3_cmp
		port map (
			clk            => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset          => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest => mm_interconnect_1_dma_rd_3_s0_waitrequest,                  --    s0.waitrequest
			s0_burstcount  => mm_interconnect_1_dma_rd_3_s0_burstcount,                   --      .burstcount
			s0_writedata   => mm_interconnect_1_dma_rd_3_s0_writedata,                    --      .writedata
			s0_address     => mm_interconnect_1_dma_rd_3_s0_address,                      --      .address
			s0_write       => mm_interconnect_1_dma_rd_3_s0_write,                        --      .write
			s0_byteenable  => mm_interconnect_1_dma_rd_3_s0_byteenable,                   --      .byteenable
			m0_waitrequest => rd_dma_3_waitrequest,                                       --    m0.waitrequest
			m0_burstcount  => rd_dma_3_burstcount,                                        --      .burstcount
			m0_writedata   => rd_dma_3_writedata,                                         --      .writedata
			m0_address     => rd_dma_3_address,                                           --      .address
			m0_write       => rd_dma_3_write,                                             --      .write
			m0_byteenable  => rd_dma_3_byteenable                                         --      .byteenable
		);

	dma_wr_0 : component PCIE_HIP_FDAS_mm_rd_transparent_0_cmp
		port map (
			clk              => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset            => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest   => mm_interconnect_0_dma_wr_0_s0_waitrequest,                  --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_dma_wr_0_s0_readdata,                     --      .readdata
			s0_readdatavalid => mm_interconnect_0_dma_wr_0_s0_readdatavalid,                --      .readdatavalid
			s0_response      => mm_interconnect_0_dma_wr_0_s0_response,                     --      .response
			s0_burstcount    => mm_interconnect_0_dma_wr_0_s0_burstcount,                   --      .burstcount
			s0_address       => mm_interconnect_0_dma_wr_0_s0_address,                      --      .address
			s0_read          => mm_interconnect_0_dma_wr_0_s0_read,                         --      .read
			m0_waitrequest   => wr_dma_0_waitrequest,                                       --    m0.waitrequest
			m0_readdata      => wr_dma_0_readdata,                                          --      .readdata
			m0_readdatavalid => wr_dma_0_readdatavalid,                                     --      .readdatavalid
			m0_response      => wr_dma_0_response,                                          --      .response
			m0_burstcount    => wr_dma_0_burstcount,                                        --      .burstcount
			m0_address       => wr_dma_0_address,                                           --      .address
			m0_read          => wr_dma_0_read                                               --      .read
		);

	dma_wr_1 : component PCIE_HIP_FDAS_mm_rd_transparent_1_cmp
		port map (
			clk              => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset            => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest   => mm_interconnect_0_dma_wr_1_s0_waitrequest,                  --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_dma_wr_1_s0_readdata,                     --      .readdata
			s0_readdatavalid => mm_interconnect_0_dma_wr_1_s0_readdatavalid,                --      .readdatavalid
			s0_response      => mm_interconnect_0_dma_wr_1_s0_response,                     --      .response
			s0_burstcount    => mm_interconnect_0_dma_wr_1_s0_burstcount,                   --      .burstcount
			s0_address       => mm_interconnect_0_dma_wr_1_s0_address,                      --      .address
			s0_read          => mm_interconnect_0_dma_wr_1_s0_read,                         --      .read
			m0_waitrequest   => wr_dma_1_waitrequest,                                       --    m0.waitrequest
			m0_readdata      => wr_dma_1_readdata,                                          --      .readdata
			m0_readdatavalid => wr_dma_1_readdatavalid,                                     --      .readdatavalid
			m0_response      => wr_dma_1_response,                                          --      .response
			m0_burstcount    => wr_dma_1_burstcount,                                        --      .burstcount
			m0_address       => wr_dma_1_address,                                           --      .address
			m0_read          => wr_dma_1_read                                               --      .read
		);

	dma_wr_2 : component PCIE_HIP_FDAS_mm_rd_transparent_2_cmp
		port map (
			clk              => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset            => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest   => mm_interconnect_0_dma_wr_2_s0_waitrequest,                  --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_dma_wr_2_s0_readdata,                     --      .readdata
			s0_readdatavalid => mm_interconnect_0_dma_wr_2_s0_readdatavalid,                --      .readdatavalid
			s0_response      => mm_interconnect_0_dma_wr_2_s0_response,                     --      .response
			s0_burstcount    => mm_interconnect_0_dma_wr_2_s0_burstcount,                   --      .burstcount
			s0_address       => mm_interconnect_0_dma_wr_2_s0_address,                      --      .address
			s0_read          => mm_interconnect_0_dma_wr_2_s0_read,                         --      .read
			m0_waitrequest   => wr_dma_2_waitrequest,                                       --    m0.waitrequest
			m0_readdata      => wr_dma_2_readdata,                                          --      .readdata
			m0_readdatavalid => wr_dma_2_readdatavalid,                                     --      .readdatavalid
			m0_response      => wr_dma_2_response,                                          --      .response
			m0_burstcount    => wr_dma_2_burstcount,                                        --      .burstcount
			m0_address       => wr_dma_2_address,                                           --      .address
			m0_read          => wr_dma_2_read                                               --      .read
		);

	dma_wr_3 : component PCIE_HIP_FDAS_mm_rd_transparent_3_cmp
		port map (
			clk              => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset            => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest   => mm_interconnect_0_dma_wr_3_s0_waitrequest,                  --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_dma_wr_3_s0_readdata,                     --      .readdata
			s0_readdatavalid => mm_interconnect_0_dma_wr_3_s0_readdatavalid,                --      .readdatavalid
			s0_response      => mm_interconnect_0_dma_wr_3_s0_response,                     --      .response
			s0_burstcount    => mm_interconnect_0_dma_wr_3_s0_burstcount,                   --      .burstcount
			s0_address       => mm_interconnect_0_dma_wr_3_s0_address,                      --      .address
			s0_read          => mm_interconnect_0_dma_wr_3_s0_read,                         --      .read
			m0_waitrequest   => wr_dma_3_waitrequest,                                       --    m0.waitrequest
			m0_readdata      => wr_dma_3_readdata,                                          --      .readdata
			m0_readdatavalid => wr_dma_3_readdatavalid,                                     --      .readdatavalid
			m0_response      => wr_dma_3_response,                                          --      .response
			m0_burstcount    => wr_dma_3_burstcount,                                        --      .burstcount
			m0_address       => wr_dma_3_address,                                           --      .address
			m0_read          => wr_dma_3_read                                               --      .read
		);

	intel_pcie_ptile_mcdma_0 : component PCIE_HIP_FDAS_intel_pcie_ptile_mcdma_0_cmp
		port map (
			app_clk                     => intel_pcie_ptile_mcdma_0_app_clk_clk,                         --           app_clk.clk
			app_rst_n                   => intel_pcie_ptile_mcdma_0_app_nreset_status_reset,             -- app_nreset_status.reset_n
			rx_pio_waitrequest_i        => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_waitrequest,        --  p0_rx_pio_master.waitrequest
			rx_pio_address_o            => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_address,            --                  .address
			rx_pio_byteenable_o         => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_byteenable,         --                  .byteenable
			rx_pio_read_o               => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_read,               --                  .read
			rx_pio_readdata_i           => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdata,           --                  .readdata
			rx_pio_readdatavalid_i      => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdatavalid,      --                  .readdatavalid
			rx_pio_write_o              => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_write,              --                  .write
			rx_pio_writedata_o          => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writedata,          --                  .writedata
			rx_pio_burstcount_o         => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_burstcount,         --                  .burstcount
			rx_pio_response_i           => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_response,           --                  .response
			rx_pio_writeresponsevalid_i => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writeresponsevalid, --                  .writeresponsevalid
			d2hdm_waitrequest_i         => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_waitrequest,         --   p0_d2hdm_master.waitrequest
			d2hdm_read_o                => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_read,                --                  .read
			d2hdm_address_o             => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_address,             --                  .address
			d2hdm_burstcount_o          => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_burstcount,          --                  .burstcount
			d2hdm_byteenable_o          => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_byteenable,          --                  .byteenable
			d2hdm_readdatavalid_i       => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdatavalid,       --                  .readdatavalid
			d2hdm_readdata_i            => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdata,            --                  .readdata
			d2hdm_response_i            => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_response,            --                  .response
			h2ddm_waitrequest_i         => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_waitrequest,         --   p0_h2ddm_master.waitrequest
			h2ddm_write_o               => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_write,               --                  .write
			h2ddm_address_o             => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_address,             --                  .address
			h2ddm_burstcount_o          => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_burstcount,          --                  .burstcount
			h2ddm_byteenable_o          => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_byteenable,          --                  .byteenable
			h2ddm_writedata_o           => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_writedata,           --                  .writedata
			usr_event_msix_valid_i      => intel_pcie_ptile_mcdma_0_p0_usr_msix_valid,                   --       p0_usr_msix.valid
			usr_event_msix_ready_o      => intel_pcie_ptile_mcdma_0_p0_usr_msix_ready,                   --                  .ready
			usr_event_msix_data_i       => intel_pcie_ptile_mcdma_0_p0_usr_msix_data,                    --                  .data
			usr_hip_tl_cfg_func_o       => open,                                                         --  p0_usr_config_tl.tl_cfg_func
			usr_hip_tl_cfg_add_o        => open,                                                         --                  .tl_cfg_add
			usr_hip_tl_cfg_ctl_o        => open,                                                         --                  .tl_cfg_ctl
			p0_link_up_o                => open,                                                         --     p0_hip_status.link_up
			p0_dl_up_o                  => open,                                                         --                  .dl_up
			p0_surprise_down_err_o      => open,                                                         --                  .surprise_down_err
			p0_ltssm_state_o            => open,                                                         --                  .ltssmstate
			refclk0                     => intel_pcie_ptile_mcdma_0_refclk0_clk,                         --           refclk0.clk
			refclk1                     => intel_pcie_ptile_mcdma_0_refclk1_clk,                         --           refclk1.clk
			ninit_done                  => intel_pcie_ptile_mcdma_0_ninit_done_reset,                    --        ninit_done.reset
			rx_n_in0                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in0,                 --        hip_serial.rx_n_in0
			rx_n_in1                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in1,                 --                  .rx_n_in1
			rx_n_in2                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in2,                 --                  .rx_n_in2
			rx_n_in3                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in3,                 --                  .rx_n_in3
			rx_n_in4                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in4,                 --                  .rx_n_in4
			rx_n_in5                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in5,                 --                  .rx_n_in5
			rx_n_in6                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in6,                 --                  .rx_n_in6
			rx_n_in7                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in7,                 --                  .rx_n_in7
			rx_n_in8                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in8,                 --                  .rx_n_in8
			rx_n_in9                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in9,                 --                  .rx_n_in9
			rx_n_in10                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in10,                --                  .rx_n_in10
			rx_n_in11                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in11,                --                  .rx_n_in11
			rx_n_in12                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in12,                --                  .rx_n_in12
			rx_n_in13                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in13,                --                  .rx_n_in13
			rx_n_in14                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in14,                --                  .rx_n_in14
			rx_n_in15                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_n_in15,                --                  .rx_n_in15
			rx_p_in0                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in0,                 --                  .rx_p_in0
			rx_p_in1                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in1,                 --                  .rx_p_in1
			rx_p_in2                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in2,                 --                  .rx_p_in2
			rx_p_in3                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in3,                 --                  .rx_p_in3
			rx_p_in4                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in4,                 --                  .rx_p_in4
			rx_p_in5                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in5,                 --                  .rx_p_in5
			rx_p_in6                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in6,                 --                  .rx_p_in6
			rx_p_in7                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in7,                 --                  .rx_p_in7
			rx_p_in8                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in8,                 --                  .rx_p_in8
			rx_p_in9                    => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in9,                 --                  .rx_p_in9
			rx_p_in10                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in10,                --                  .rx_p_in10
			rx_p_in11                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in11,                --                  .rx_p_in11
			rx_p_in12                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in12,                --                  .rx_p_in12
			rx_p_in13                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in13,                --                  .rx_p_in13
			rx_p_in14                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in14,                --                  .rx_p_in14
			rx_p_in15                   => intel_pcie_ptile_mcdma_0_hip_serial_rx_p_in15,                --                  .rx_p_in15
			tx_n_out0                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out0,                --                  .tx_n_out0
			tx_n_out1                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out1,                --                  .tx_n_out1
			tx_n_out2                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out2,                --                  .tx_n_out2
			tx_n_out3                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out3,                --                  .tx_n_out3
			tx_n_out4                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out4,                --                  .tx_n_out4
			tx_n_out5                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out5,                --                  .tx_n_out5
			tx_n_out6                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out6,                --                  .tx_n_out6
			tx_n_out7                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out7,                --                  .tx_n_out7
			tx_n_out8                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out8,                --                  .tx_n_out8
			tx_n_out9                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out9,                --                  .tx_n_out9
			tx_n_out10                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out10,               --                  .tx_n_out10
			tx_n_out11                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out11,               --                  .tx_n_out11
			tx_n_out12                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out12,               --                  .tx_n_out12
			tx_n_out13                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out13,               --                  .tx_n_out13
			tx_n_out14                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out14,               --                  .tx_n_out14
			tx_n_out15                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_n_out15,               --                  .tx_n_out15
			tx_p_out0                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out0,                --                  .tx_p_out0
			tx_p_out1                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out1,                --                  .tx_p_out1
			tx_p_out2                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out2,                --                  .tx_p_out2
			tx_p_out3                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out3,                --                  .tx_p_out3
			tx_p_out4                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out4,                --                  .tx_p_out4
			tx_p_out5                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out5,                --                  .tx_p_out5
			tx_p_out6                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out6,                --                  .tx_p_out6
			tx_p_out7                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out7,                --                  .tx_p_out7
			tx_p_out8                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out8,                --                  .tx_p_out8
			tx_p_out9                   => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out9,                --                  .tx_p_out9
			tx_p_out10                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out10,               --                  .tx_p_out10
			tx_p_out11                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out11,               --                  .tx_p_out11
			tx_p_out12                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out12,               --                  .tx_p_out12
			tx_p_out13                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out13,               --                  .tx_p_out13
			tx_p_out14                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out14,               --                  .tx_p_out14
			tx_p_out15                  => intel_pcie_ptile_mcdma_0_hip_serial_tx_p_out15,               --                  .tx_p_out15
			pin_perst_n                 => intel_pcie_ptile_mcdma_0_pin_perst_reset_n                    --         pin_perst.reset_n
		);

	reset_bridge_0 : component PCIE_HIP_FDAS_reset_bridge_0_cmp
		port map (
			clk         => intel_pcie_ptile_mcdma_0_app_clk_clk,             --       clk.clk
			in_reset_n  => intel_pcie_ptile_mcdma_0_app_nreset_status_reset, --  in_reset.reset_n
			out_reset_n => reset_out_reset_n                                 -- out_reset.reset_n
		);

	rxm_bar2_0 : component PCIE_HIP_FDAS_mm_transparent_no_burst_pio_0_cmp
		port map (
			clk                   => intel_pcie_ptile_mcdma_0_app_clk_clk,                       -- clock.clk
			reset                 => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- reset.reset
			s0_waitrequest        => mm_interconnect_2_rxm_bar2_0_s0_waitrequest,                --    s0.waitrequest
			s0_readdata           => mm_interconnect_2_rxm_bar2_0_s0_readdata,                   --      .readdata
			s0_readdatavalid      => mm_interconnect_2_rxm_bar2_0_s0_readdatavalid,              --      .readdatavalid
			s0_writeresponsevalid => mm_interconnect_2_rxm_bar2_0_s0_writeresponsevalid,         --      .writeresponsevalid
			s0_response           => mm_interconnect_2_rxm_bar2_0_s0_response,                   --      .response
			s0_writedata          => mm_interconnect_2_rxm_bar2_0_s0_writedata,                  --      .writedata
			s0_address            => mm_interconnect_2_rxm_bar2_0_s0_address,                    --      .address
			s0_write              => mm_interconnect_2_rxm_bar2_0_s0_write,                      --      .write
			s0_read               => mm_interconnect_2_rxm_bar2_0_s0_read,                       --      .read
			s0_byteenable         => mm_interconnect_2_rxm_bar2_0_s0_byteenable,                 --      .byteenable
			m0_waitrequest        => rxm_bar2_0_m0_waitrequest,                                  --    m0.waitrequest
			m0_readdata           => rxm_bar2_0_m0_readdata,                                     --      .readdata
			m0_readdatavalid      => rxm_bar2_0_m0_readdatavalid,                                --      .readdatavalid
			m0_writeresponsevalid => rxm_bar2_0_m0_writeresponsevalid,                           --      .writeresponsevalid
			m0_response           => rxm_bar2_0_m0_response,                                     --      .response
			m0_writedata          => rxm_bar2_0_m0_writedata,                                    --      .writedata
			m0_address            => rxm_bar2_0_m0_address,                                      --      .address
			m0_write              => rxm_bar2_0_m0_write,                                        --      .write
			m0_read               => rxm_bar2_0_m0_read,                                         --      .read
			m0_byteenable         => rxm_bar2_0_m0_byteenable                                    --      .byteenable
		);

	mm_interconnect_0 : component PCIE_HIP_FDAS_altera_mm_interconnect_1920_yasd64i_cmp
		port map (
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_address                                      => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_address,           --                                        intel_pcie_ptile_mcdma_0_p0_d2hdm_master.address
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_waitrequest                                  => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_waitrequest,       --                                                                                .waitrequest
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_burstcount                                   => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_burstcount,        --                                                                                .burstcount
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_byteenable                                   => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_byteenable,        --                                                                                .byteenable
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_read                                         => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_read,              --                                                                                .read
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdata                                     => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdata,          --                                                                                .readdata
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdatavalid                                => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_readdatavalid,     --                                                                                .readdatavalid
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_response                                     => intel_pcie_ptile_mcdma_0_p0_d2hdm_master_response,          --                                                                                .response
			dma_wr_0_s0_address                                                                   => mm_interconnect_0_dma_wr_0_s0_address,                      --                                                                     dma_wr_0_s0.address
			dma_wr_0_s0_read                                                                      => mm_interconnect_0_dma_wr_0_s0_read,                         --                                                                                .read
			dma_wr_0_s0_readdata                                                                  => mm_interconnect_0_dma_wr_0_s0_readdata,                     --                                                                                .readdata
			dma_wr_0_s0_burstcount                                                                => mm_interconnect_0_dma_wr_0_s0_burstcount,                   --                                                                                .burstcount
			dma_wr_0_s0_readdatavalid                                                             => mm_interconnect_0_dma_wr_0_s0_readdatavalid,                --                                                                                .readdatavalid
			dma_wr_0_s0_waitrequest                                                               => mm_interconnect_0_dma_wr_0_s0_waitrequest,                  --                                                                                .waitrequest
			dma_wr_0_s0_response                                                                  => mm_interconnect_0_dma_wr_0_s0_response,                     --                                                                                .response
			dma_wr_1_s0_address                                                                   => mm_interconnect_0_dma_wr_1_s0_address,                      --                                                                     dma_wr_1_s0.address
			dma_wr_1_s0_read                                                                      => mm_interconnect_0_dma_wr_1_s0_read,                         --                                                                                .read
			dma_wr_1_s0_readdata                                                                  => mm_interconnect_0_dma_wr_1_s0_readdata,                     --                                                                                .readdata
			dma_wr_1_s0_burstcount                                                                => mm_interconnect_0_dma_wr_1_s0_burstcount,                   --                                                                                .burstcount
			dma_wr_1_s0_readdatavalid                                                             => mm_interconnect_0_dma_wr_1_s0_readdatavalid,                --                                                                                .readdatavalid
			dma_wr_1_s0_waitrequest                                                               => mm_interconnect_0_dma_wr_1_s0_waitrequest,                  --                                                                                .waitrequest
			dma_wr_1_s0_response                                                                  => mm_interconnect_0_dma_wr_1_s0_response,                     --                                                                                .response
			dma_wr_2_s0_address                                                                   => mm_interconnect_0_dma_wr_2_s0_address,                      --                                                                     dma_wr_2_s0.address
			dma_wr_2_s0_read                                                                      => mm_interconnect_0_dma_wr_2_s0_read,                         --                                                                                .read
			dma_wr_2_s0_readdata                                                                  => mm_interconnect_0_dma_wr_2_s0_readdata,                     --                                                                                .readdata
			dma_wr_2_s0_burstcount                                                                => mm_interconnect_0_dma_wr_2_s0_burstcount,                   --                                                                                .burstcount
			dma_wr_2_s0_readdatavalid                                                             => mm_interconnect_0_dma_wr_2_s0_readdatavalid,                --                                                                                .readdatavalid
			dma_wr_2_s0_waitrequest                                                               => mm_interconnect_0_dma_wr_2_s0_waitrequest,                  --                                                                                .waitrequest
			dma_wr_2_s0_response                                                                  => mm_interconnect_0_dma_wr_2_s0_response,                     --                                                                                .response
			dma_wr_3_s0_address                                                                   => mm_interconnect_0_dma_wr_3_s0_address,                      --                                                                     dma_wr_3_s0.address
			dma_wr_3_s0_read                                                                      => mm_interconnect_0_dma_wr_3_s0_read,                         --                                                                                .read
			dma_wr_3_s0_readdata                                                                  => mm_interconnect_0_dma_wr_3_s0_readdata,                     --                                                                                .readdata
			dma_wr_3_s0_burstcount                                                                => mm_interconnect_0_dma_wr_3_s0_burstcount,                   --                                                                                .burstcount
			dma_wr_3_s0_readdatavalid                                                             => mm_interconnect_0_dma_wr_3_s0_readdatavalid,                --                                                                                .readdatavalid
			dma_wr_3_s0_waitrequest                                                               => mm_interconnect_0_dma_wr_3_s0_waitrequest,                  --                                                                                .waitrequest
			dma_wr_3_s0_response                                                                  => mm_interconnect_0_dma_wr_3_s0_response,                     --                                                                                .response
			dma_wr_0_reset_reset_bridge_in_reset_reset                                            => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, --                                            dma_wr_0_reset_reset_bridge_in_reset.reset
			intel_pcie_ptile_mcdma_0_p0_d2hdm_master_translator_reset_reset_bridge_in_reset_reset => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- intel_pcie_ptile_mcdma_0_p0_d2hdm_master_translator_reset_reset_bridge_in_reset.reset
			intel_pcie_ptile_mcdma_0_app_clk_clk                                                  => intel_pcie_ptile_mcdma_0_app_clk_clk                        --                                                intel_pcie_ptile_mcdma_0_app_clk.clk
		);

	mm_interconnect_1 : component PCIE_HIP_FDAS_altera_mm_interconnect_1920_j3desai_cmp
		port map (
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_address                                      => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_address,           --                                        intel_pcie_ptile_mcdma_0_p0_h2ddm_master.address
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_waitrequest                                  => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_waitrequest,       --                                                                                .waitrequest
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_burstcount                                   => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_burstcount,        --                                                                                .burstcount
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_byteenable                                   => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_byteenable,        --                                                                                .byteenable
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_write                                        => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_write,             --                                                                                .write
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_writedata                                    => intel_pcie_ptile_mcdma_0_p0_h2ddm_master_writedata,         --                                                                                .writedata
			dma_rd_0_s0_address                                                                   => mm_interconnect_1_dma_rd_0_s0_address,                      --                                                                     dma_rd_0_s0.address
			dma_rd_0_s0_write                                                                     => mm_interconnect_1_dma_rd_0_s0_write,                        --                                                                                .write
			dma_rd_0_s0_writedata                                                                 => mm_interconnect_1_dma_rd_0_s0_writedata,                    --                                                                                .writedata
			dma_rd_0_s0_burstcount                                                                => mm_interconnect_1_dma_rd_0_s0_burstcount,                   --                                                                                .burstcount
			dma_rd_0_s0_byteenable                                                                => mm_interconnect_1_dma_rd_0_s0_byteenable,                   --                                                                                .byteenable
			dma_rd_0_s0_waitrequest                                                               => mm_interconnect_1_dma_rd_0_s0_waitrequest,                  --                                                                                .waitrequest
			dma_rd_1_s0_address                                                                   => mm_interconnect_1_dma_rd_1_s0_address,                      --                                                                     dma_rd_1_s0.address
			dma_rd_1_s0_write                                                                     => mm_interconnect_1_dma_rd_1_s0_write,                        --                                                                                .write
			dma_rd_1_s0_writedata                                                                 => mm_interconnect_1_dma_rd_1_s0_writedata,                    --                                                                                .writedata
			dma_rd_1_s0_burstcount                                                                => mm_interconnect_1_dma_rd_1_s0_burstcount,                   --                                                                                .burstcount
			dma_rd_1_s0_byteenable                                                                => mm_interconnect_1_dma_rd_1_s0_byteenable,                   --                                                                                .byteenable
			dma_rd_1_s0_waitrequest                                                               => mm_interconnect_1_dma_rd_1_s0_waitrequest,                  --                                                                                .waitrequest
			dma_rd_2_s0_address                                                                   => mm_interconnect_1_dma_rd_2_s0_address,                      --                                                                     dma_rd_2_s0.address
			dma_rd_2_s0_write                                                                     => mm_interconnect_1_dma_rd_2_s0_write,                        --                                                                                .write
			dma_rd_2_s0_writedata                                                                 => mm_interconnect_1_dma_rd_2_s0_writedata,                    --                                                                                .writedata
			dma_rd_2_s0_burstcount                                                                => mm_interconnect_1_dma_rd_2_s0_burstcount,                   --                                                                                .burstcount
			dma_rd_2_s0_byteenable                                                                => mm_interconnect_1_dma_rd_2_s0_byteenable,                   --                                                                                .byteenable
			dma_rd_2_s0_waitrequest                                                               => mm_interconnect_1_dma_rd_2_s0_waitrequest,                  --                                                                                .waitrequest
			dma_rd_3_s0_address                                                                   => mm_interconnect_1_dma_rd_3_s0_address,                      --                                                                     dma_rd_3_s0.address
			dma_rd_3_s0_write                                                                     => mm_interconnect_1_dma_rd_3_s0_write,                        --                                                                                .write
			dma_rd_3_s0_writedata                                                                 => mm_interconnect_1_dma_rd_3_s0_writedata,                    --                                                                                .writedata
			dma_rd_3_s0_burstcount                                                                => mm_interconnect_1_dma_rd_3_s0_burstcount,                   --                                                                                .burstcount
			dma_rd_3_s0_byteenable                                                                => mm_interconnect_1_dma_rd_3_s0_byteenable,                   --                                                                                .byteenable
			dma_rd_3_s0_waitrequest                                                               => mm_interconnect_1_dma_rd_3_s0_waitrequest,                  --                                                                                .waitrequest
			dma_rd_0_reset_reset_bridge_in_reset_reset                                            => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, --                                            dma_rd_0_reset_reset_bridge_in_reset.reset
			intel_pcie_ptile_mcdma_0_p0_h2ddm_master_translator_reset_reset_bridge_in_reset_reset => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv, -- intel_pcie_ptile_mcdma_0_p0_h2ddm_master_translator_reset_reset_bridge_in_reset.reset
			intel_pcie_ptile_mcdma_0_app_clk_clk                                                  => intel_pcie_ptile_mcdma_0_app_clk_clk                        --                                                intel_pcie_ptile_mcdma_0_app_clk.clk
		);

	mm_interconnect_2 : component PCIE_HIP_FDAS_altera_mm_interconnect_1920_jrv6pua_cmp
		port map (
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_address                                      => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_address,            --                                        intel_pcie_ptile_mcdma_0_p0_rx_pio_master.address
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_waitrequest                                  => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_waitrequest,        --                                                                                 .waitrequest
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_burstcount                                   => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_burstcount,         --                                                                                 .burstcount
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_byteenable                                   => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_byteenable,         --                                                                                 .byteenable
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_read                                         => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_read,               --                                                                                 .read
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdata                                     => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdata,           --                                                                                 .readdata
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdatavalid                                => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_readdatavalid,      --                                                                                 .readdatavalid
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_write                                        => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_write,              --                                                                                 .write
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writedata                                    => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writedata,          --                                                                                 .writedata
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_response                                     => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_response,           --                                                                                 .response
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writeresponsevalid                           => intel_pcie_ptile_mcdma_0_p0_rx_pio_master_writeresponsevalid, --                                                                                 .writeresponsevalid
			rxm_bar2_0_s0_address                                                                  => mm_interconnect_2_rxm_bar2_0_s0_address,                      --                                                                    rxm_bar2_0_s0.address
			rxm_bar2_0_s0_write                                                                    => mm_interconnect_2_rxm_bar2_0_s0_write,                        --                                                                                 .write
			rxm_bar2_0_s0_read                                                                     => mm_interconnect_2_rxm_bar2_0_s0_read,                         --                                                                                 .read
			rxm_bar2_0_s0_readdata                                                                 => mm_interconnect_2_rxm_bar2_0_s0_readdata,                     --                                                                                 .readdata
			rxm_bar2_0_s0_writedata                                                                => mm_interconnect_2_rxm_bar2_0_s0_writedata,                    --                                                                                 .writedata
			rxm_bar2_0_s0_byteenable                                                               => mm_interconnect_2_rxm_bar2_0_s0_byteenable,                   --                                                                                 .byteenable
			rxm_bar2_0_s0_readdatavalid                                                            => mm_interconnect_2_rxm_bar2_0_s0_readdatavalid,                --                                                                                 .readdatavalid
			rxm_bar2_0_s0_waitrequest                                                              => mm_interconnect_2_rxm_bar2_0_s0_waitrequest,                  --                                                                                 .waitrequest
			rxm_bar2_0_s0_response                                                                 => mm_interconnect_2_rxm_bar2_0_s0_response,                     --                                                                                 .response
			rxm_bar2_0_s0_writeresponsevalid                                                       => mm_interconnect_2_rxm_bar2_0_s0_writeresponsevalid,           --                                                                                 .writeresponsevalid
			rxm_bar2_0_reset_reset_bridge_in_reset_reset                                           => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv,   --                                           rxm_bar2_0_reset_reset_bridge_in_reset.reset
			intel_pcie_ptile_mcdma_0_p0_rx_pio_master_translator_reset_reset_bridge_in_reset_reset => intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv,   -- intel_pcie_ptile_mcdma_0_p0_rx_pio_master_translator_reset_reset_bridge_in_reset.reset
			intel_pcie_ptile_mcdma_0_app_clk_clk                                                   => intel_pcie_ptile_mcdma_0_app_clk_clk                          --                                                 intel_pcie_ptile_mcdma_0_app_clk.clk
		);

	intel_pcie_ptile_mcdma_0_app_nreset_status_reset_ports_inv <= not intel_pcie_ptile_mcdma_0_app_nreset_status_reset;

end architecture rtl; -- of PCIE_HIP_FDAS
