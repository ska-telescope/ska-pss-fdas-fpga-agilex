----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2023 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
--
-- VHDL Architecture conv_lib.conv.scm
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 18:31:57 11/09/2023
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

LIBRARY conv_lib;

ARCHITECTURE scm OF conv IS

  -- Architecture declarations
  type word32_array_t is array (natural range <>) of std_logic_vector(31 downto 0);

  -- Internal signal declarations
  SIGNAL ready2_s                 : std_logic;                                                  --       .sink_ready
  SIGNAL mcdataout2_s             : std_logic_vector(ifft_g*32-1 DOWNTO 0);
  SIGNAL mcdataout1_s             : std_logic_vector(31 DOWNTO 0);
  SIGNAL coef_mcrden_s            : std_logic_vector(ifft_g*ifft_loop_g-1 DOWNTO 0);
  SIGNAL coef_mcwren_s            : std_logic_vector(ifft_g*ifft_loop_g-1 DOWNTO 0);
  SIGNAL coef_rdaddrout_s         : std_logic_vector(9 DOWNTO 0);
  SIGNAL coef_rdenout_s           : std_logic_vector(ifft_loop_g-1 DOWNTO 0);
  SIGNAL data5_s                  : word32_array_t(2*ifft_g-1 DOWNTO 0);
  SIGNAL data6_s                  : word32_array_t(2*ifft_g*ifft_loop_g DOWNTO 0);
  SIGNAL data5_0_s                : std_logic_vector(31 DOWNTO 0);
  SIGNAL loop_addr5_s             : std_logic_vector(ifft_loop_bits_g-1 DOWNTO 0);
  SIGNAL done6_0_s                : std_logic;
  SIGNAL eof1_s                   : std_logic;
  SIGNAL eof2_s                   : std_logic;
  SIGNAL eof3_s                   : std_logic;
  SIGNAL eof4_s                   : std_logic_vector(2*ifft_g-1 DOWNTO 0);
  SIGNAL idata1_s                 : std_logic_vector(31 DOWNTO 0);
  SIGNAL idata2_s                 : std_logic_vector(31 DOWNTO 0);
  SIGNAL data3_s                  : cmplx_array_t(2*ifft_g-1 DOWNTO 0);
  SIGNAL coefconj_s               : cmplx_array_t(ifft_g-1 DOWNTO 0);
  SIGNAL coef_s                   : cmplx_array_t(ifft_g-1 DOWNTO 0);
  SIGNAL rdata1_s                 : std_logic_vector(31 DOWNTO 0);
  SIGNAL rdata2_s                 : std_logic_vector(31 DOWNTO 0);                              -- az
  SIGNAL data4_s                  : cmplx_array_t(2*ifft_g-1 DOWNTO 0);
  SIGNAL ready1_s                 : std_logic;
  SIGNAL loop_addr2_s             : std_logic_vector(ifft_loop_bits_g-1 DOWNTO 0);
  SIGNAL sof1_s                   : std_logic;
  SIGNAL sof2_s                   : std_logic;
  SIGNAL sof3_s                   : std_logic;
  SIGNAL sof4_s                   : std_logic_vector(2*ifft_g-1 DOWNTO 0);
  SIGNAL valid1_s                 : std_logic;
  SIGNAL valid2_s                 : std_logic;
  SIGNAL valid3_s                 : std_logic;
  SIGNAL valid4_s                 : std_logic_vector(2*ifft_g-1 DOWNTO 0);
  SIGNAL valid5_0_s               : std_logic;
  SIGNAL clken_s                  : std_logic;
  SIGNAL rden_s                   : std_logic_vector(2*ifft_g*ifft_loop_g DOWNTO 0);
  SIGNAL rddata_s                 : std_logic_vector((2*ifft_g*ifft_loop_g+1)*32-1 DOWNTO 0);
  SIGNAL rdaddr0_s                : std_logic_vector(abits_g-1 DOWNTO 0);
  SIGNAL rdaddr_s                 : std_logic_vector(abits_g-1 DOWNTO 0);
  SIGNAL sof5_0_s                 : std_logic;
  SIGNAL eof5_0_s                 : std_logic;
  SIGNAL rdeof_s                  : std_logic;
  SIGNAL valid5_s                 : std_logic;
  SIGNAL sof5_s                   : std_logic;
  SIGNAL eof5_s                   : std_logic;
  SIGNAL wren5_s                  : std_logic_vector(ifft_loop_g-1 DOWNTO 0);
  SIGNAL ctrl3_s                  : std_logic_vector(ifft_loop_bits_g+1 DOWNTO 0);
  SIGNAL loop_addr3_s             : std_logic_vector(ifft_loop_bits_g-1 DOWNTO 0);
  SIGNAL ctrl2_s                  : std_logic_vector(ifft_loop_bits_g+1 DOWNTO 0);
  SIGNAL filter_coefficients_s    : filter_coefficients_out_t;
  SIGNAL filter_coefficients_rd_s : std_logic_vector(31 DOWNTO 0);
  SIGNAL fft_results_s            : fft_results_out_t;
  SIGNAL valid_0_s                : std_logic;
  SIGNAL overflow_s               : std_logic_vector(2*ifft_g*ifft_loop_g DOWNTO 0);
  SIGNAL ready6_s                 : std_logic_vector(2*ifft_g*ifft_loop_g DOWNTO 0);
  SIGNAL avail6_s                 : std_logic_vector(2*ifft_g*ifft_loop_g DOWNTO 0);
  SIGNAL avail_s                  : std_logic;
  SIGNAL ready3_0_s               : std_logic;
  SIGNAL readye_s                 : std_logic_vector(ifft_loop_g-1 DOWNTO 0);
  SIGNAL overflow_lat_s           : std_logic_vector(84 DOWNTO 0);
  SIGNAL row0_delay_s             : std_logic_vector(9 DOWNTO 0);
  SIGNAL rst_sys_n_d1             : std_logic;
  SIGNAL tie1_s                   : std_logic;
  SIGNAL rst_sys_1_n_s            : std_logic;
  SIGNAL rst_sys_0_n_s            : std_logic;


  -- Component Declarations
  COMPONENT conv_coef_str
  GENERIC (
    dbits_g : natural;
    depth_g : natural;
    abits_g : natural;
    loop_g  : natural
  );
  PORT (
    CLK_SYS      : IN     std_logic ;
    RST_SYS_N    : IN     std_logic ;
    RDATAOUT     : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    IDATACONJOUT : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    RDATACONJOUT : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    IDATAOUT     : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    RDEN         : IN     std_logic_vector (loop_g-1 DOWNTO 0);
    RDADDR       : IN     std_logic_vector (abits_g-1 DOWNTO 0);
    CLK_MC       : IN     std_logic ;
    RST_MC_N     : IN     std_logic ;
    MCADDR       : IN     std_logic_vector (abits_g DOWNTO 0);
    MCRDEN       : IN     std_logic_vector (loop_g-1 DOWNTO 0);
    MCDATAOUT    : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    MCWREN       : IN     std_logic_vector (loop_g-1 DOWNTO 0);
    MCDATA       : IN     std_logic_vector (dbits_g-1 DOWNTO 0)
  );
  END COMPONENT conv_coef_str;
  COMPONENT conv_fft
  GENERIC (
    ptsnum_g : natural
  );
  PORT (
    CLK_SYS   : IN     std_logic ;
    RST_SYS_N : IN     std_logic ;
    READY     : IN     std_logic ;
    RDATA     : IN     std_logic_vector (31 DOWNTO 0);
    IDATA     : IN     std_logic_vector (31 DOWNTO 0);
    VALID     : IN     std_logic ;
    SOF       : IN     std_logic ;
    EOF       : IN     std_logic ;
    RDATAOUT  : OUT    std_logic_vector (31 DOWNTO 0);
    IDATAOUT  : OUT    std_logic_vector (31 DOWNTO 0);
    VALIDOUT  : OUT    std_logic ;
    SOFOUT    : OUT    std_logic ;
    EOFOUT    : OUT    std_logic ;
    READYOUT  : OUT    std_logic ;
    SYNC      : IN     std_logic 
  );
  END COMPONENT conv_fft;
  COMPONENT conv_fft_str
  GENERIC (
    dbits_g     : natural;
    depth_g     : natural;
    abits_g     : natural;
    pages_g     : natural;    -- lte 2**pgbits_g
    pgbits_g    : natural;
    loop_g      : natural;    -- number of output frame repeats lte 2**loop_bits_g 
    loop_bits_g : natural
  );
  PORT (
    CLK_SYS        : IN     std_logic ;
    RST_SYS_N      : IN     std_logic ;
    RDATAOUT       : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    IDATAOUT       : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    VALIDOUT       : OUT    std_logic ;
    SOFOUT         : OUT    std_logic ;
    EOFOUT         : OUT    std_logic ;
    LOOP_ADDROUT   : OUT    std_logic_vector (loop_bits_g-1 DOWNTO 0);
    READYOUT       : OUT    std_logic ;
    COEF_RDENOUT   : OUT    std_logic_vector (loop_g-1 DOWNTO 0);
    COEF_RDADDROUT : OUT    std_logic_vector (abits_g-1 DOWNTO 0);
    RDATA          : IN     std_logic_vector (dbits_g-1 DOWNTO 0);
    IDATA          : IN     std_logic_vector (dbits_g-1 DOWNTO 0);
    VALID          : IN     std_logic ;
    SOF            : IN     std_logic ;
    EOF            : IN     std_logic ;
    LOOP_NUM       : IN     std_logic_vector (loop_bits_g DOWNTO 0);
    CONV_ENABLE    : IN     std_logic ;
    SYNC           : IN     std_logic ;
    READY          : IN     std_logic_vector (loop_g-1 DOWNTO 0);
    CLK_MC         : IN     std_logic ;
    RST_MC_N       : IN     std_logic ;
    MCADDR         : IN     std_logic_vector (abits_g DOWNTO 0);
    MCRDEN         : IN     std_logic ;
    MCDATAOUT      : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    DONEOUT        : OUT    std_logic ;
    OVERFLOW       : OUT    std_logic 
  );
  END COMPONENT conv_fft_str;
  COMPONENT conv_ifft
  GENERIC (
    ptsnum_g : natural
  );
  PORT (
    CLK_SYS   : IN     std_logic ;
    RST_SYS_N : IN     std_logic ;
    RDATAOUT  : OUT    std_logic_vector (31 DOWNTO 0);
    IDATAOUT  : OUT    std_logic_vector (31 DOWNTO 0);
    VALIDOUT  : OUT    std_logic ;
    SOFOUT    : OUT    std_logic ;
    EOFOUT    : OUT    std_logic ;
    RDATA     : IN     std_logic_vector (31 DOWNTO 0);
    IDATA     : IN     std_logic_vector (31 DOWNTO 0);
    VALID     : IN     std_logic ;
    SOF       : IN     std_logic ;
    EOF       : IN     std_logic ;
    SYNC      : IN     std_logic 
  );
  END COMPONENT conv_ifft;
  COMPONENT conv_ifft_ctrl
  GENERIC (
    stages_g    : natural;
    loop_g      : natural;    --lte 2**loop_bits_g
    loop_bits_g : natural
  );
  PORT (
    SOF          : IN     std_logic ;
    EOF          : IN     std_logic ;
    VALID        : IN     std_logic ;
    READY        : IN     std_logic ;
    SYNC         : IN     std_logic ;
    LOOP_NUM     : IN     std_logic_vector (loop_bits_g DOWNTO 0);
    CLK          : IN     std_logic ;
    CLKEN        : IN     std_logic ;
    RST_N        : IN     std_logic ;
    SOFOUT       : OUT    std_logic ;
    EOFOUT       : OUT    std_logic ;
    VALIDOUT     : OUT    std_logic ;
    LOOP_ADDROUT : OUT    std_logic_vector (loop_bits_g-1 DOWNTO 0);
    WRENOUT      : OUT    std_logic_vector (loop_g-1 DOWNTO 0)
  );
  END COMPONENT conv_ifft_ctrl;
  COMPONENT conv_mult
  PORT (
    CLK_SYS      : IN     std_logic ;
    ICOEF        : IN     std_logic_vector (31 DOWNTO 0);
    ICOEFCONJ    : IN     std_logic_vector (31 DOWNTO 0);
    IDATA        : IN     std_logic_vector (31 DOWNTO 0);
    RCOEF        : IN     std_logic_vector (31 DOWNTO 0);
    RCOEFCONJ    : IN     std_logic_vector (31 DOWNTO 0);
    RDATA        : IN     std_logic_vector (31 DOWNTO 0);
    RST_SYS_N    : IN     std_logic ;
    VALID        : IN     std_logic ;
    IDATACONJOUT : OUT    std_logic_vector (31 DOWNTO 0); -- result
    IDATAOUT     : OUT    std_logic_vector (31 DOWNTO 0);
    RDATACONJOUT : OUT    std_logic_vector (31 DOWNTO 0); -- result
    RDATAOUT     : OUT    std_logic_vector (31 DOWNTO 0)
  );
  END COMPONENT conv_mult;
  COMPONENT conv_pwr
  PORT (
    CLK_SYS   : IN     std_logic ;
    EOF       : IN     std_logic ;
    IDATA     : IN     std_logic_vector (31 DOWNTO 0); -- az
    RDATA     : IN     std_logic_vector (31 DOWNTO 0);
    RST_SYS_N : IN     std_logic ;
    SOF       : IN     std_logic ;
    SYNC      : IN     std_logic ;
    VALID     : IN     std_logic ;
    DATAOUT   : OUT    std_logic_vector (31 DOWNTO 0);
    EOFOUT    : OUT    std_logic ;
    SOFOUT    : OUT    std_logic ;
    VALIDOUT  : OUT    std_logic 
  );
  END COMPONENT conv_pwr;
  COMPONENT conv_result_str
  GENERIC (
    dbits_g  : natural;
    depth_g  : natural;
    abits_g  : natural;
    pages_g  : natural;    -- lte 2**pgbits_g
    pgbits_g : natural
  );
  PORT (
    CLK_SYS   : IN     std_logic ;
    RST_SYS_N : IN     std_logic ;
    RDADDR    : IN     std_logic_vector (abits_g-1 DOWNTO 0);
    RDEN      : IN     std_logic ;
    RDEOF     : IN     std_logic ;
    DATAOUT   : OUT    std_logic_vector (dbits_g-1 DOWNTO 0);
    DATA      : IN     std_logic_vector (dbits_g-1 DOWNTO 0);
    VALID     : IN     std_logic ;
    SOF       : IN     std_logic ;
    EOF       : IN     std_logic ;
    SYNC      : IN     std_logic ;
    AVAILOUT  : OUT    std_logic ;
    READYOUT  : OUT    std_logic ;
    OVERFLOW  : OUT    std_logic ;
    DONEOUT   : OUT    std_logic 
  );
  END COMPONENT conv_result_str;
  COMPONENT convmci
  PORT (
    MCADDR                 : IN     std_logic_vector (19 DOWNTO 0);
    MCDATAIN               : IN     std_logic_vector (31 DOWNTO 0);
    MCDATAOUT              : OUT    std_logic_vector (31 DOWNTO 0);
    MCRWN                  : IN     std_logic ;
    MCMS                   : IN     std_logic ;
    CLK_MC                 : IN     std_logic ;
    RST_MC_N               : IN     std_logic ;
    FILTER_COEFFICIENTS    : OUT    filter_coefficients_out_t ;
    FILTER_COEFFICIENTS_RD : IN     std_logic_vector (31 DOWNTO 0);
    FFT_RESULTS            : OUT    fft_results_out_t ;
    FFT_RESULTS_RD         : IN     std_logic_vector (31 DOWNTO 0);
    ROW0_DELAY             : OUT    std_logic_vector (9 DOWNTO 0);
    OVERFLOW               : IN     std_logic_vector (84 DOWNTO 0)
  );
  END COMPONENT convmci;
  COMPONENT convreset_sync
  PORT (
    RST_N       : IN     std_logic ;
    CLK         : IN     std_logic ;
    RST_OUT_0_N : OUT    std_logic ;
    RST_OUT_1_N : OUT    std_logic 
  );
  END COMPONENT convreset_sync;
  COMPONENT fop_str
  GENERIC (
    ddr_g            : natural;
    abits_g          : natural;
    ifft_g           : natural;
    ifft_loop_g      : natural;    -- number of output frame repeats lte 2**ifft_loop_bits_g
    ifft_loop_bits_g : natural;
    fop_num_bits_g   : natural;
    delay_g          : natural;
    delaybits_g      : natural
  );
  PORT (
    CLK_SYS       : IN     std_logic ;
    RST_SYS_N     : IN     std_logic ;
    RDADDROUT     : OUT    std_logic_vector (abits_g-1 DOWNTO 0);
    RDADDR0OUT    : OUT    std_logic_vector (abits_g-1 DOWNTO 0);
    RDENOUT       : OUT    std_logic_vector (2*ifft_g*ifft_loop_g DOWNTO 0);
    RDEOFOUT      : OUT    std_logic ;
    RDDATA        : IN     std_logic_vector ((2*ifft_g*ifft_loop_g+1)*32-1 DOWNTO 0);
    DDR_WAITREQ   : IN     std_logic ;
    AVAIL         : IN     std_logic ;
    DDR_ADDROUT   : OUT    std_logic_vector (25 DOWNTO 0);
    DDR_DATAOUT   : OUT    std_logic_vector (ddr_g*512-1 DOWNTO 0);
    DDR_VALIDOUT  : OUT    std_logic ;
    DONEOUT       : OUT    std_logic ;
    CONV_DONEOUT  : OUT    std_logic ;
    IFFT_LOOP_NUM : IN     std_logic_vector (ifft_loop_bits_g DOWNTO 0);
    FOP_NUM       : IN     std_logic_vector (fop_num_bits_g-1 DOWNTO 0);
    OVERLAP_SIZE  : IN     std_logic_vector (abits_g-1 DOWNTO 0);
    ROW0_DELAY    : IN     std_logic_vector (abits_g-1 DOWNTO 0);
    PAGE_START    : IN     std_logic_vector (25 DOWNTO 0);
    SYNC          : IN     std_logic ;
    CONV_ENABLE   : IN     std_logic 
  );
  END COMPONENT fop_str;
  COMPONENT retime
  GENERIC (
    dataw_g  : natural;
    stages_g : natural
  );
  PORT (
    DATA    : IN     std_logic_vector (dataw_g-1 DOWNTO 0);
    DE      : IN     std_logic ;
    SYNC    : IN     std_logic ;
    CLK     : IN     std_logic ;
    CLKEN   : IN     std_logic ;
    RST_N   : IN     std_logic ;
    DATAOUT : OUT    std_logic_vector (dataw_g-1 DOWNTO 0);
    DEOUT   : OUT    std_logic 
  );
  END COMPONENT retime;

  -- Optional embedded configurations
  -- pragma synthesis_off
  FOR ALL : conv_fft USE ENTITY conv_lib.conv_fft;
  FOR ALL : conv_fft_str USE ENTITY conv_lib.conv_fft_str;
  FOR ALL : conv_ifft_ctrl USE ENTITY conv_lib.conv_ifft_ctrl;
  FOR pwr1_i : conv_pwr USE ENTITY conv_lib.conv_pwr;
  FOR result_str0_i : conv_result_str USE ENTITY conv_lib.conv_result_str;
  FOR ALL : convmci USE ENTITY conv_lib.convmci;
  FOR ALL : convreset_sync USE ENTITY conv_lib.convreset_sync;
  FOR ALL : fop_str USE ENTITY conv_lib.fop_str;
  FOR ALL : retime USE ENTITY conv_lib.retime;
  -- pragma synthesis_on


BEGIN
  -- Architecture concurrent statements
  -- HDL Embedded Text Block 1 eb1
  -- eb1 1
  decode_mcen_filt: for f in 0 to ifft_g-1 generate
    decode_mcen_rpt:  for r in 0 to ifft_loop_g-1 generate
      coef_mcrden_s(f*ifft_loop_g+r) <= filter_coefficients_s.rden when to_integer(unsigned(filter_coefficients_s.addr(16 downto 11))) = r*ifft_g+f else
                                   '0';
      coef_mcwren_s(f*ifft_loop_g+r) <= filter_coefficients_s.wren when to_integer(unsigned(filter_coefficients_s.addr(16 downto 11))) = r*ifft_g+f else
                                   '0';
    end generate decode_mcen_rpt;
  end generate decode_mcen_filt;
  
  
  
  

  -- HDL Embedded Text Block 2 eb2
  -- eb2 2
  loop_addr3_s <= ctrl3_s(ifft_loop_bits_g+1 downto 2);
  sof3_s <= ctrl3_s(0);
  eof3_s <= ctrl3_s(1);
                                          

  -- HDL Embedded Text Block 3 eb3
  -- eb3 3
  ctrl2_s <= loop_addr2_s & eof2_s & sof2_s;                                        

  -- HDL Embedded Text Block 4 eb4
  -- eb4 4
  valid_0_s <= VALID and ready1_s;
  READYOUT <= ready1_s;
  tie1_s <= '1';                               

  -- HDL Embedded Text Block 5 eb5
  -- eb5 5
  clken_s <= '1';
  ready3_0_s <= '1';                                        

  -- HDL Embedded Text Block 6 eb6
  -- eb6 6
  genrddata: for i in 0 to 2*ifft_g*ifft_loop_g generate
    rddata_s((i+1)*32-1 downto i*32) <= data6_s(i);
  end generate;                                        

  -- HDL Embedded Text Block 7 eb7
  -- eb7 7
  -- or mcdataout from conv_coef_str modules
  gen_coef_mcdataout : process (mcdataout2_s)
    variable mcdataout_v : std_logic_vector(31 downto 0);
  begin
    mcdataout_v := (others => '0');
    for i in 0 to ifft_g-1 loop
      mcdataout_v := mcdataout_v or mcdataout2_s((i+1)*32-1 downto i*32);
    end loop;
    filter_coefficients_rd_s <= mcdataout_v;
  end process gen_coef_mcdataout;                                       
  
  

  -- HDL Embedded Text Block 8 eb8
  -- eb8 8
  avail_s <= avail6_s(2*ifft_g*to_integer(unsigned(IFFT_LOOP_NUM)));                                        

  -- HDL Embedded Text Block 9 eb9
  -- eb9 9
  -- extract ready for each repeat
  extract_ready: for r in 0 to ifft_loop_g-1 generate
    readye_s(r) <= ready6_s(2*ifft_g*(r+1));
  end generate extract_ready;

  -- HDL Embedded Text Block 10 eb10
  -- eb10 10
  --------------------------------------------------------------------------
  -- latch overflow alarms
  --------------------------------------------------------------------------
  latch_alarms : process (CLK_SYS,rst_sys_0_n_s)
  begin
    if rst_sys_0_n_s='0' then
      overflow_lat_s <= (others => '0');
    elsif rising_edge(CLK_SYS) then
      -- on trigger shift clear latched overflow alarms
      if CONV_TRIGGER='1' then
        overflow_lat_s <= (others => '0');
      end if;
      -- latch overflow indicators
      for i in 0 to 2*ifft_g*ifft_loop_g loop
        if overflow_s(i)='1' then
          overflow_lat_s(i) <= '1';
        end if;
      end loop;
    end if;
  end process latch_alarms;
                                          


  -- Instance port mappings.
  fft_i : conv_fft
    GENERIC MAP (
      ptsnum_g => fft_g
    )
    PORT MAP (
      CLK_SYS   => CLK_SYS,
      RST_SYS_N => rst_sys_0_n_s,
      READY     => ready2_s,
      RDATA     => RDATA,
      IDATA     => IDATA,
      VALID     => VALID,
      SOF       => SOF,
      EOF       => EOF,
      RDATAOUT  => rdata1_s,
      IDATAOUT  => idata1_s,
      VALIDOUT  => valid1_s,
      SOFOUT    => sof1_s,
      EOFOUT    => eof1_s,
      READYOUT  => ready1_s,
      SYNC      => CONV_TRIGGER
    );
  fft_str_i : conv_fft_str
    GENERIC MAP (
      dbits_g     => 32,
      depth_g     => fft_g,
      abits_g     => abits_g,
      pages_g     => 4,                -- lte 2**pgbits_g
      pgbits_g    => 2,
      loop_g      => ifft_loop_g,      -- number of output frame repeats lte 2**loop_bits_g 
      loop_bits_g => ifft_loop_bits_g
    )
    PORT MAP (
      CLK_SYS => CLK_SYS,
      RST_SYS_N => rst_sys_0_n_s,
      RDATAOUT => rdata2_s,
      IDATAOUT => idata2_s,
      VALIDOUT => valid2_s,
      SOFOUT => sof2_s,
      EOFOUT => eof2_s,
      LOOP_ADDROUT => loop_addr2_s,
      READYOUT => ready2_s,
      COEF_RDENOUT => coef_rdenout_s,
      COEF_RDADDROUT => coef_rdaddrout_s,
      RDATA => rdata1_s,
      IDATA => idata1_s,
      VALID => valid1_s,
      SOF => sof1_s,
      EOF => eof1_s,
      LOOP_NUM => IFFT_LOOP_NUM,
      CONV_ENABLE => CONV_ENABLE,
      SYNC => CONV_TRIGGER,
      READY => readye_s,
      CLK_MC => CLK_MC,
      RST_MC_N => RST_MC_N,
      MCDATAOUT => mcdataout1_s,
      DONEOUT => MCREADYOUT,
      MCADDR => fft_results_s.addr,
      MCRDEN => fft_results_s.rden,
      OVERFLOW => open
    );
  ifft_ctrl_i : conv_ifft_ctrl
    GENERIC MAP (
      stages_g    => 4,
      loop_g      => ifft_loop_g,      --lte 2**loop_bits_g
      loop_bits_g => ifft_loop_bits_g
    )
    PORT MAP (
      SOF          => sof4_s(0),
      EOF          => eof4_s(0),
      VALID        => valid4_s(0),
      READY        => tie1_s,
      SYNC         => CONV_TRIGGER,
      LOOP_NUM     => IFFT_LOOP_NUM,
      CLK          => CLK_SYS,
      CLKEN        => clken_s,
      RST_N        => rst_sys_0_n_s,
      SOFOUT       => sof5_s,
      EOFOUT       => eof5_s,
      VALIDOUT     => valid5_s,
      LOOP_ADDROUT => loop_addr5_s,
      WRENOUT      => wren5_s
    );
  pwr1_i : conv_pwr
    PORT MAP (
      CLK_SYS   => CLK_SYS,
      EOF       => EOF,
      IDATA     => IDATA,
      RDATA     => RDATA,
      RST_SYS_N => rst_sys_1_n_s,
      SOF       => SOF,
      SYNC      => CONV_TRIGGER,
      VALID     => valid_0_s,
      DATAOUT   => data5_0_s,
      EOFOUT    => eof5_0_s,
      SOFOUT    => sof5_0_s,
      VALIDOUT  => valid5_0_s
    );
  result_str0_i : conv_result_str
    GENERIC MAP (
      dbits_g  => 32,
      depth_g  => fft_g,
      abits_g  => abits_g,
      pages_g  => res_pages_g+4,      -- lte 2**pgbits_g
      pgbits_g => integer(ceil(log2(real(res_pages_g+4))))
    )
    PORT MAP (
      CLK_SYS   => CLK_SYS,
      RST_SYS_N => rst_sys_1_n_s,
      RDADDR    => rdaddr0_s,
      RDEN      => rden_s(0),
      RDEOF     => rdeof_s,
      DATAOUT   => data6_s(0),
      DATA      => data5_0_s,
      VALID     => valid5_0_s,
      SOF       => sof5_0_s,
      EOF       => eof5_0_s,
      SYNC      => CONV_TRIGGER,
      AVAILOUT  => avail6_s(0),
      READYOUT  => ready6_s(0),
      OVERFLOW  => overflow_s(0),
      DONEOUT   => done6_0_s
    );
  mci_i : convmci
    PORT MAP (
      MCADDR                 => MCADDR,
      MCDATAIN               => MCDATA,
      MCDATAOUT              => MCDATAOUT,
      MCRWN                  => MCRWN,
      MCMS                   => MCMS,
      CLK_MC                 => CLK_MC,
      RST_MC_N               => RST_MC_N,
      FILTER_COEFFICIENTS    => filter_coefficients_s,
      FILTER_COEFFICIENTS_RD => filter_coefficients_rd_s,
      FFT_RESULTS            => fft_results_s,
      FFT_RESULTS_RD         => mcdataout1_s,
      ROW0_DELAY             => row0_delay_s,
      OVERFLOW               => overflow_lat_s
    );
  convreset_i : convreset_sync
    PORT MAP (
      RST_N       => RST_SYS_N,
      CLK         => CLK_SYS,
      RST_OUT_0_N => rst_sys_0_n_s,
      RST_OUT_1_N => rst_sys_1_n_s
    );
  fop_str_i : fop_str
    GENERIC MAP (
      ddr_g            => ddr_g,
      abits_g          => abits_g,
      ifft_g           => ifft_g,
      ifft_loop_g      => ifft_loop_g,      -- number of output frame repeats lte 2**ifft_loop_bits_g
      ifft_loop_bits_g => ifft_loop_bits_g,
      fop_num_bits_g   => fop_num_bits_g,
      delay_g          => 2,
      delaybits_g      => 3
    )
    PORT MAP (
      CLK_SYS => CLK_SYS,
      RST_SYS_N => rst_sys_1_n_s,
      RDADDROUT => rdaddr_s,
      RDADDR0OUT => rdaddr0_s,
      RDENOUT => rden_s,
      RDEOFOUT => rdeof_s,
      RDDATA => rddata_s,
      DDR_WAITREQ => DDR_WAITREQ,
      AVAIL => avail_s,
      DDR_ADDROUT => DDR_ADDROUT,
      DDR_DATAOUT => DDR_DATAOUT,
      DDR_VALIDOUT => DDR_VALIDOUT,
      DONEOUT => SEGDONEOUT,
      CONV_DONEOUT => CONV_DONEOUT,
      IFFT_LOOP_NUM => IFFT_LOOP_NUM,
      FOP_NUM => FOP_NUM,
      OVERLAP_SIZE => OVERLAP_SIZE,
      ROW0_DELAY => row0_delay_s,
      PAGE_START => PAGE_START,
      SYNC => CONV_TRIGGER,
      CONV_ENABLE => CONV_ENABLE
    );
  retime1_i : retime
    GENERIC MAP (
      dataw_g  => ifft_loop_bits_g+2,
      stages_g => 5
    )
    PORT MAP (
      DATA    => ctrl2_s,
      DE      => valid2_s,
      SYNC    => CONV_TRIGGER,
      CLK     => CLK_SYS,
      CLKEN   => clken_s,
      RST_N   => rst_sys_1_n_s,
      DATAOUT => ctrl3_s,
      DEOUT   => valid3_s
    );

  g0: FOR i IN 0 TO ifft_g-1 GENERATE
  -- Optional embedded configurations
  -- pragma synthesis_off
  FOR ALL : conv_coef_str USE ENTITY conv_lib.conv_coef_str;
  FOR ALL : conv_mult USE ENTITY conv_lib.conv_mult;
  -- pragma synthesis_on

  BEGIN
    coef_i : conv_coef_str
      GENERIC MAP (
        dbits_g => 32,
        depth_g => fft_g,
        abits_g => abits_g,
        loop_g  => ifft_loop_g
      )
      PORT MAP (
        CLK_SYS => CLK_SYS,
        RST_SYS_N => rst_sys_1_n_s,
        RDEN => coef_rdenout_s,
        RDADDR => coef_rdaddrout_s,
        CLK_MC => CLK_MC,
        RST_MC_N => RST_MC_N,
        RDATAOUT => coef_s(i).RE,
        IDATACONJOUT => coefconj_s(i).IM,
        RDATACONJOUT => coefconj_s(i).RE,
        IDATAOUT => coef_s(i).IM,
        MCADDR => filter_coefficients_s.addr(abits_g downto 0),
        MCRDEN => coef_mcrden_s((i+1)*ifft_loop_g-1 downto i*ifft_loop_g),
        MCDATAOUT => mcdataout2_s((i+1)*32-1 downto i*32),
        MCWREN => coef_mcwren_s((i+1)*ifft_loop_g-1 downto i*ifft_loop_g),
        MCDATA => filter_coefficients_s.wr
      );
    mult_i : conv_mult
      PORT MAP (
        CLK_SYS => CLK_SYS,
        IDATA => idata2_s,
        RDATA => rdata2_s,
        RST_SYS_N => rst_sys_0_n_s,
        VALID => valid2_s,
        ICOEF => coef_s(i).IM,
        ICOEFCONJ => coefconj_s(i).IM,
        RCOEF => coef_s(i).RE,
        RCOEFCONJ => coefconj_s(i).RE,
        IDATACONJOUT => data3_s(2*i+1).IM,
        IDATAOUT => data3_s(2*i).IM,
        RDATACONJOUT => data3_s(2*i+1).RE,
        RDATAOUT => data3_s(2*i).RE
      );
  END GENERATE g0;

  g1: FOR i IN 0 TO 2*ifft_g-1 GENERATE
  -- Optional embedded configurations
  -- pragma synthesis_off
  FOR ALL : conv_ifft USE ENTITY conv_lib.conv_ifft;
  FOR pwr_i : conv_pwr USE ENTITY conv_lib.conv_pwr;
  -- pragma synthesis_on

  BEGIN
    pwr_i : conv_pwr
      PORT MAP (
        CLK_SYS => CLK_SYS,
        RST_SYS_N => rst_sys_0_n_s,
        EOF => eof4_s(i),
        IDATA => data4_s(i).IM,
        RDATA => data4_s(i).RE,
        SOF => sof4_s(i),
        SYNC => '0',
        VALID => valid4_s(i),
        DATAOUT => data5_s(i),
        EOFOUT => open,
        SOFOUT => open,
        VALIDOUT => open
      );
    ifft_i : conv_ifft
      GENERIC MAP (
        ptsnum_g => fft_g
      )
      PORT MAP (
        CLK_SYS => CLK_SYS,
        RST_SYS_N => rst_sys_1_n_s,
        VALID => valid3_s,
        SOF => sof3_s,
        EOF => eof3_s,
        SYNC => CONV_TRIGGER,
        RDATAOUT => data4_s(i).RE,
        IDATAOUT => data4_s(i).IM,
        VALIDOUT => valid4_s(i),
        SOFOUT => sof4_s(i),
        EOFOUT => eof4_s(i),
        RDATA => data3_s(i).RE,
        IDATA => data3_s(i).IM
      );
  END GENERATE g1;

  g2: FOR r IN 0 TO ifft_loop_g-1 GENERATE
  BEGIN
    g3: FOR f IN 0 TO 2*ifft_g-1 GENERATE
    -- Optional embedded configurations
    -- pragma synthesis_off
    FOR result_str_i : conv_result_str USE ENTITY conv_lib.conv_result_str;
    -- pragma synthesis_on

    BEGIN
      result_str_i : conv_result_str
        GENERIC MAP (
          dbits_g  => 32,
          depth_g  => fft_g,
          abits_g  => abits_g,
          pages_g  => res_pages_g,          -- lte 2**pgbits_g
          pgbits_g => integer(ceil(log2(real(res_pages_g))))
        )
        PORT MAP (
          CLK_SYS => CLK_SYS,
          RST_SYS_N => rst_sys_1_n_s,
          RDADDR => rdaddr_s,
          RDEOF => rdeof_s,
          SOF => sof5_s,
          EOF => eof5_s,
          SYNC => CONV_TRIGGER,
          RDEN => rden_s(r*2*ifft_g+f+1),
          DATAOUT => data6_s(r*2*ifft_g+f+1),
          DATA => data5_s(f),
          VALID => wren5_s(r),
          AVAILOUT => avail6_s(r*2*ifft_g+f+1),
          READYOUT => ready6_s(r*2*ifft_g+f+1),
          OVERFLOW => overflow_s(r*2*ifft_g+f+1),
          DONEOUT => open
        );
    END GENERATE g3;

  END GENERATE g2;

END ARCHITECTURE scm;
