----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.conv_fft.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 12:05:04 18/07/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library conv_lib;
library fft1024;

entity conv_fft is
  generic( 
    ptsnum_g : natural
  );
  port( 
    CLK_SYS   : in     std_logic;
    RST_SYS_N : in     std_logic;
    READY     : in     std_logic;
    RDATA     : in     std_logic_vector (31 downto 0);
    IDATA     : in     std_logic_vector (31 downto 0);
    VALID     : in     std_logic;
    SOF       : in     std_logic;
    EOF       : in     std_logic;
    RDATAOUT  : out    std_logic_vector (31 downto 0);
    IDATAOUT  : out    std_logic_vector (31 downto 0);
    VALIDOUT  : out    std_logic;
    SOFOUT    : out    std_logic;
    EOFOUT    : out    std_logic;
    READYOUT  : out    std_logic;
    SYNC      : in     std_logic
  );

-- Declarations

end entity conv_fft ;

