----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity cld_lib.cld.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 13:26:50 13/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY cld IS
  GENERIC( 
    ddr_g                    : integer;    --number of DDR Interfaces
    fft_ddr_addr_num_g       : integer;    --Number of DDR locations to read for an FFT
    fop_ddr_addr_max_width_g : integer;    --Number of counter bits to support the address for reading of the FOP from DDR memory
    fft_ddr_addr_num_width_g : integer;    --Number of counter bits to support ddr_addr_num_g
    fft_g                    : integer;    --Number of samples in an FFT
    fft_count_width_g        : integer;    --Number of counter bits  to support fft_g
    sample_count_width_g     : integer;    --Number of counter bits to support fop_g
    fifo_waddr_width_g       : integer;    --Number of counter bits to support write locations
    fifo_raddr_width_g       : integer     --Number of counter bits to support read locations
  );
  PORT( 
    cld_enable     : IN     std_logic;
    cld_page       : IN     std_logic_vector (31 DOWNTO 0);
    cld_trigger    : IN     std_logic;
    clk_sys        : IN     std_logic;
    data_valid     : IN     std_logic;
    ddr_data       : IN     std_logic_vector (512*ddr_g -1  DOWNTO 0);
    fop_sample_num : IN     std_logic_vector (22 DOWNTO 0);
    overlap_int    : IN     std_logic_vector (4 DOWNTO 0);
    overlap_rem    : IN     std_logic_vector (4 DOWNTO 0);
    overlap_size   : IN     std_logic_vector (9  DOWNTO 0);
    ready          : IN     std_logic;
    rst_sys_n      : IN     std_logic;
    wait_request   : IN     std_logic;
    cld_done       : OUT    std_logic;
    conv_data      : OUT    std_logic_vector (63  DOWNTO 0);
    conv_req       : OUT    std_logic;
    ddr_addr       : OUT    std_logic_vector (31 DOWNTO 0);
    ddr_read       : OUT    std_logic;
    eof            : OUT    std_logic;
    fft_sample     : OUT    std_logic_vector (9  DOWNTO 0);
    sof            : OUT    std_logic;
    valid          : OUT    std_logic
  );

-- Declarations

END ENTITY cld ;

