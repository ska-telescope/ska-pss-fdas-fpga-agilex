-- ifft1024.vhd

-- Generated using ACDS version 22.2 94

library IEEE;
library intel_FPGA_unified_fft_103;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ifft1024 is
	port (
		clk        : in  std_logic                     := '0';             --    clk.clk
		rst        : in  std_logic                     := '0';             --    rst.reset_n
		validIn    : in  std_logic_vector(0 downto 0)  := (others => '0'); --   sink.valid
		channelIn  : in  std_logic_vector(7 downto 0)  := (others => '0'); --       .channel
		d          : in  std_logic_vector(63 downto 0) := (others => '0'); --       .data
		validOut   : out std_logic_vector(0 downto 0);                     -- source.valid
		channelOut : out std_logic_vector(7 downto 0);                     --       .channel
		q          : out std_logic_vector(63 downto 0)                     --       .data
	);
end entity ifft1024;

architecture rtl of ifft1024 is
	component ifft1024_intel_FPGA_unified_fft_103_ua3wp3i_cmp is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst            : in  std_logic                     := 'X';             -- reset_n
			validIn        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			channelIn      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			in_d_real_tpl  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_d_imag_tpl  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			validOut       : out std_logic_vector(0 downto 0);                     -- valid
			channelOut     : out std_logic_vector(7 downto 0);                     -- channel
			out_q_real_tpl : out std_logic_vector(31 downto 0);                    -- data
			out_q_imag_tpl : out std_logic_vector(31 downto 0)                     -- data
		);
	end component ifft1024_intel_FPGA_unified_fft_103_ua3wp3i_cmp;

	signal intel_fpga_unified_fft_0_out_q_imag_tpl : std_logic_vector(31 downto 0); -- port fragment
	signal intel_fpga_unified_fft_0_out_q_real_tpl : std_logic_vector(31 downto 0); -- port fragment

	for intel_fpga_unified_fft_0 : ifft1024_intel_FPGA_unified_fft_103_ua3wp3i_cmp
		use entity intel_FPGA_unified_fft_103.ifft1024_intel_FPGA_unified_fft_103_ua3wp3i;
begin

	intel_fpga_unified_fft_0 : component ifft1024_intel_FPGA_unified_fft_103_ua3wp3i_cmp
		port map (
			clk                         => clk,                                                  --    clk.clk
			rst                         => rst,                                                  --    rst.reset_n
			validIn                     => validIn,                                              --   sink.valid
			channelIn                   => channelIn,                                            --       .channel
			in_d_imag_tpl(31 downto 0)  => d(63 downto 32),                                      --       .data
			in_d_real_tpl(31 downto 0)  => d(31 downto 0),                                       --       .data
			validOut                    => validOut,                                             -- source.valid
			channelOut                  => channelOut,                                           --       .channel
			out_q_imag_tpl(31 downto 0) => intel_fpga_unified_fft_0_out_q_imag_tpl(31 downto 0), --       .data
			out_q_real_tpl(31 downto 0) => intel_fpga_unified_fft_0_out_q_real_tpl(31 downto 0)  --       .data
		);

	q <= intel_FPGA_unified_fft_0_out_q_imag_tpl(31 downto 0) & intel_FPGA_unified_fft_0_out_q_real_tpl(31 downto 0);

end architecture rtl; -- of ifft1024
