----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity ctrl_lib.ctrl_func.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 11:59:37 17/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ctrl_func is
  port( 
    cld_done           : in     std_logic;
    clk_sys            : in     std_logic;
    conv_done          : in     std_logic;
    conv_waitreq       : in     std_logic;
    conv_wr_en         : in     std_logic;
    dm_trig            : in     std_logic;
    hsum_done          : in     std_logic;
    hsum_rd_en         : in     std_logic;
    hsum_valid         : in     std_logic;
    hsum_waitreq       : in     std_logic;
    man_cld_en         : in     std_logic;
    man_cld_pause_cnt  : in     std_logic_vector (31 downto 0);
    man_cld_pause_en   : in     std_logic;
    man_cld_pause_rst  : in     std_logic;
    man_cld_trig       : in     std_logic;
    man_conv_en        : in     std_logic;
    man_conv_pause_cnt : in     std_logic_vector (31 downto 0);
    man_conv_pause_en  : in     std_logic;
    man_conv_pause_rst : in     std_logic;
    man_conv_trig      : in     std_logic;
    man_hsum_en        : in     std_logic;
    man_hsum_pause_cnt : in     std_logic_vector (31 downto 0);
    man_hsum_pause_en  : in     std_logic;
    man_hsum_pause_rst : in     std_logic;
    man_hsum_trig      : in     std_logic;
    man_override       : in     std_logic;
    page               : in     std_logic;
    rst_sys_n          : in     std_logic;
    cld_enable         : out    std_logic;
    cld_page           : out    std_logic_vector (31 downto 0);
    cld_paused         : out    std_logic;
    cld_proc_time      : out    std_logic_vector (31 downto 0);
    cld_trigger        : out    std_logic;
    conv_enable        : out    std_logic;
    conv_page          : out    std_logic_vector (31 downto 0);
    conv_paused        : out    std_logic;
    conv_proc_time     : out    std_logic_vector (31 downto 0);
    conv_req_cnt       : out    std_logic_vector (31 downto 0);
    conv_trigger       : out    std_logic;
    hsum_enable        : out    std_logic;
    hsum_page          : out    std_logic_vector (31 downto 0);
    hsum_paused        : out    std_logic;
    hsum_proc_time     : out    std_logic_vector (31 downto 0);
    hsum_rec_cnt       : out    std_logic_vector (31 downto 0);
    hsum_req_cnt       : out    std_logic_vector (31 downto 0);
    hsum_trigger       : out    std_logic;
    latched_cld_done   : out    std_logic;
    latched_conv_done  : out    std_logic;
    latched_hsum_done  : out    std_logic
  );

-- Declarations

end entity ctrl_func ;

