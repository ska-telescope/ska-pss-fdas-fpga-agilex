-- ed_sim.vhd

-- Generated using ACDS version 22.2 94

library IEEE;
library ed_sim_emif_cal;
library ed_sim_emif_fm_0;
library ed_sim_local_reset_combiner;
library ed_sim_local_reset_source;
library ed_sim_mem;
library ed_sim_ninit_done;
library ed_sim_pll_ref_clk_source;
library ed_sim_sim_checker;
library ed_sim_tg;
library altera_mm_interconnect_1920;
library altera_reset_controller_1921;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ed_sim is
	port (
		sim_checker_traffic_gen_pass         : out std_logic;  --        sim_checker.traffic_gen_pass
		sim_checker_traffic_gen_fail         : out std_logic;  --                   .traffic_gen_fail
		sim_checker_traffic_gen_timeout      : out std_logic;  --                   .traffic_gen_timeout
		cal_status_checker_local_cal_success : out std_logic;  -- cal_status_checker.local_cal_success
		cal_status_checker_local_cal_fail    : out std_logic   --                   .local_cal_fail
	);
end entity ed_sim;

architecture rtl of ed_sim is
	component ed_sim_emif_cal_cmp is
		port (
			calbus_read_0          : out std_logic;                                          -- calbus_read
			calbus_write_0         : out std_logic;                                          -- calbus_write
			calbus_address_0       : out std_logic_vector(19 downto 0);                      -- calbus_address
			calbus_wdata_0         : out std_logic_vector(31 downto 0);                      -- calbus_wdata
			calbus_rdata_0         : in  std_logic_vector(31 downto 0)   := (others => 'X'); -- calbus_rdata
			calbus_seq_param_tbl_0 : in  std_logic_vector(4095 downto 0) := (others => 'X'); -- calbus_seq_param_tbl
			calbus_clk             : out std_logic                                           -- clk
		);
	end component ed_sim_emif_cal_cmp;

	component ed_sim_emif_fm_0_cmp is
		port (
			local_reset_req      : in    std_logic                       := 'X';             -- local_reset_req
			local_reset_done     : out   std_logic;                                          -- local_reset_done
			pll_ref_clk          : in    std_logic                       := 'X';             -- clk
			pll_ref_clk_out      : out   std_logic;                                          -- clk
			pll_locked           : out   std_logic;                                          -- pll_locked
			oct_rzqin            : in    std_logic                       := 'X';             -- oct_rzqin
			mem_ck               : out   std_logic_vector(0 downto 0);                       -- mem_ck
			mem_ck_n             : out   std_logic_vector(0 downto 0);                       -- mem_ck_n
			mem_a                : out   std_logic_vector(16 downto 0);                      -- mem_a
			mem_act_n            : out   std_logic_vector(0 downto 0);                       -- mem_act_n
			mem_ba               : out   std_logic_vector(1 downto 0);                       -- mem_ba
			mem_bg               : out   std_logic_vector(1 downto 0);                       -- mem_bg
			mem_cke              : out   std_logic_vector(0 downto 0);                       -- mem_cke
			mem_cs_n             : out   std_logic_vector(0 downto 0);                       -- mem_cs_n
			mem_odt              : out   std_logic_vector(0 downto 0);                       -- mem_odt
			mem_reset_n          : out   std_logic_vector(0 downto 0);                       -- mem_reset_n
			mem_par              : out   std_logic_vector(0 downto 0);                       -- mem_par
			mem_alert_n          : in    std_logic_vector(0 downto 0)    := (others => 'X'); -- mem_alert_n
			mem_dqs              : inout std_logic_vector(8 downto 0)    := (others => 'X'); -- mem_dqs
			mem_dqs_n            : inout std_logic_vector(8 downto 0)    := (others => 'X'); -- mem_dqs_n
			mem_dq               : inout std_logic_vector(71 downto 0)   := (others => 'X'); -- mem_dq
			mem_dbi_n            : inout std_logic_vector(8 downto 0)    := (others => 'X'); -- mem_dbi_n
			local_cal_success    : out   std_logic;                                          -- local_cal_success
			local_cal_fail       : out   std_logic;                                          -- local_cal_fail
			emif_usr_reset_n     : out   std_logic;                                          -- reset_n
			emif_usr_clk         : out   std_logic;                                          -- clk
			amm_ready_0          : out   std_logic;                                          -- waitrequest_n
			amm_read_0           : in    std_logic                       := 'X';             -- read
			amm_write_0          : in    std_logic                       := 'X';             -- write
			amm_address_0        : in    std_logic_vector(26 downto 0)   := (others => 'X'); -- address
			amm_readdata_0       : out   std_logic_vector(575 downto 0);                     -- readdata
			amm_writedata_0      : in    std_logic_vector(575 downto 0)  := (others => 'X'); -- writedata
			amm_burstcount_0     : in    std_logic_vector(6 downto 0)    := (others => 'X'); -- burstcount
			amm_byteenable_0     : in    std_logic_vector(71 downto 0)   := (others => 'X'); -- byteenable
			amm_readdatavalid_0  : out   std_logic;                                          -- readdatavalid
			calbus_read          : in    std_logic                       := 'X';             -- calbus_read
			calbus_write         : in    std_logic                       := 'X';             -- calbus_write
			calbus_address       : in    std_logic_vector(19 downto 0)   := (others => 'X'); -- calbus_address
			calbus_wdata         : in    std_logic_vector(31 downto 0)   := (others => 'X'); -- calbus_wdata
			calbus_rdata         : out   std_logic_vector(31 downto 0);                      -- calbus_rdata
			calbus_seq_param_tbl : out   std_logic_vector(4095 downto 0);                    -- calbus_seq_param_tbl
			calbus_clk           : in    std_logic                       := 'X'              -- clk
		);
	end component ed_sim_emif_fm_0_cmp;

	component ed_sim_local_reset_combiner_cmp is
		port (
			local_reset_req_out_0 : out std_logic;        -- local_reset_req
			local_reset_done_in_0 : in  std_logic := 'X'; -- local_reset_done
			clk                   : in  std_logic := 'X'; -- clk
			reset_n               : in  std_logic := 'X'; -- pll_locked
			local_reset_req       : in  std_logic := 'X'; -- local_reset_req
			local_reset_done      : out std_logic         -- local_reset_done
		);
	end component ed_sim_local_reset_combiner_cmp;

	component ed_sim_local_reset_source_cmp is
		port (
			local_reset_req  : out std_logic;        -- local_reset_req
			local_reset_done : in  std_logic := 'X'  -- local_reset_done
		);
	end component ed_sim_local_reset_source_cmp;

	component ed_sim_mem_cmp is
		port (
			mem_ck      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_ck
			mem_ck_n    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_ck_n
			mem_a       : in    std_logic_vector(16 downto 0) := (others => 'X'); -- mem_a
			mem_act_n   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_act_n
			mem_ba      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_ba
			mem_bg      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_bg
			mem_cke     : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cke
			mem_cs_n    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cs_n
			mem_odt     : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_odt
			mem_reset_n : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_reset_n
			mem_par     : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_par
			mem_alert_n : out   std_logic_vector(0 downto 0);                     -- mem_alert_n
			mem_dqs     : inout std_logic_vector(8 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n   : inout std_logic_vector(8 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_dq      : inout std_logic_vector(71 downto 0) := (others => 'X'); -- mem_dq
			mem_dbi_n   : inout std_logic_vector(8 downto 0)  := (others => 'X')  -- mem_dbi_n
		);
	end component ed_sim_mem_cmp;

	component ed_sim_ninit_done_cmp is
		port (
			ninit_done : out std_logic   -- reset
		);
	end component ed_sim_ninit_done_cmp;

	component ed_sim_pll_ref_clk_source_cmp is
		generic (
			CLOCK_RATE : positive := 33333000;
			CLOCK_UNIT : positive := 1
		);
		port (
			clk : out std_logic   -- clk
		);
	end component ed_sim_pll_ref_clk_source_cmp;

	component ed_sim_sim_checker_cmp is
		port (
			traffic_gen_pass_0    : in  std_logic := 'X'; -- traffic_gen_pass
			traffic_gen_fail_0    : in  std_logic := 'X'; -- traffic_gen_fail
			traffic_gen_timeout_0 : in  std_logic := 'X'; -- traffic_gen_timeout
			traffic_gen_pass      : out std_logic;        -- traffic_gen_pass
			traffic_gen_fail      : out std_logic;        -- traffic_gen_fail
			traffic_gen_timeout   : out std_logic;        -- traffic_gen_timeout
			local_cal_success_0   : in  std_logic := 'X'; -- local_cal_success
			local_cal_fail_0      : in  std_logic := 'X'; -- local_cal_fail
			local_cal_success     : out std_logic;        -- local_cal_success
			local_cal_fail        : out std_logic         -- local_cal_fail
		);
	end component ed_sim_sim_checker_cmp;

	component ed_sim_tg_cmp is
		port (
			emif_usr_reset_n      : in  std_logic                      := 'X';             -- reset_n
			ninit_done            : in  std_logic                      := 'X';             -- reset
			emif_usr_clk          : in  std_logic                      := 'X';             -- clk
			amm_ready_0           : in  std_logic                      := 'X';             -- waitrequest_n
			amm_read_0            : out std_logic;                                         -- read
			amm_write_0           : out std_logic;                                         -- write
			amm_address_0         : out std_logic_vector(33 downto 0);                     -- address
			amm_readdata_0        : in  std_logic_vector(575 downto 0) := (others => 'X'); -- readdata
			amm_writedata_0       : out std_logic_vector(575 downto 0);                    -- writedata
			amm_burstcount_0      : out std_logic_vector(6 downto 0);                      -- burstcount
			amm_byteenable_0      : out std_logic_vector(71 downto 0);                     -- byteenable
			amm_readdatavalid_0   : in  std_logic                      := 'X';             -- readdatavalid
			traffic_gen_pass_0    : out std_logic;                                         -- traffic_gen_pass
			traffic_gen_fail_0    : out std_logic;                                         -- traffic_gen_fail
			traffic_gen_timeout_0 : out std_logic                                          -- traffic_gen_timeout
		);
	end component ed_sim_tg_cmp;

	component ed_sim_altera_mm_interconnect_1920_2l4tnfq_cmp is
		port (
			tg_ctrl_amm_0_address                                      : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- address
			tg_ctrl_amm_0_waitrequest                                  : out std_logic;                                         -- waitrequest
			tg_ctrl_amm_0_burstcount                                   : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- burstcount
			tg_ctrl_amm_0_byteenable                                   : in  std_logic_vector(71 downto 0)  := (others => 'X'); -- byteenable
			tg_ctrl_amm_0_read                                         : in  std_logic                      := 'X';             -- read
			tg_ctrl_amm_0_readdata                                     : out std_logic_vector(575 downto 0);                    -- readdata
			tg_ctrl_amm_0_readdatavalid                                : out std_logic;                                         -- readdatavalid
			tg_ctrl_amm_0_write                                        : in  std_logic                      := 'X';             -- write
			tg_ctrl_amm_0_writedata                                    : in  std_logic_vector(575 downto 0) := (others => 'X'); -- writedata
			emif_fm_0_ctrl_amm_0_address                               : out std_logic_vector(26 downto 0);                     -- address
			emif_fm_0_ctrl_amm_0_write                                 : out std_logic;                                         -- write
			emif_fm_0_ctrl_amm_0_read                                  : out std_logic;                                         -- read
			emif_fm_0_ctrl_amm_0_readdata                              : in  std_logic_vector(575 downto 0) := (others => 'X'); -- readdata
			emif_fm_0_ctrl_amm_0_writedata                             : out std_logic_vector(575 downto 0);                    -- writedata
			emif_fm_0_ctrl_amm_0_burstcount                            : out std_logic_vector(6 downto 0);                      -- burstcount
			emif_fm_0_ctrl_amm_0_byteenable                            : out std_logic_vector(71 downto 0);                     -- byteenable
			emif_fm_0_ctrl_amm_0_readdatavalid                         : in  std_logic                      := 'X';             -- readdatavalid
			emif_fm_0_ctrl_amm_0_waitrequest                           : in  std_logic                      := 'X';             -- waitrequest
			tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			emif_fm_0_emif_usr_clk_clk                                 : in  std_logic                      := 'X'              -- clk
		);
	end component ed_sim_altera_mm_interconnect_1920_2l4tnfq_cmp;

	component altera_reset_controller_cmp is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller_cmp;

	signal pll_ref_clk_source_clk_clk                                 : std_logic;                       -- pll_ref_clk_source:clk -> emif_fm_0:pll_ref_clk
	signal emif_cal_emif_calbus_clk_clk                               : std_logic;                       -- emif_cal:calbus_clk -> emif_fm_0:calbus_clk
	signal emif_fm_0_emif_usr_clk_clk                                 : std_logic;                       -- emif_fm_0:emif_usr_clk -> [mm_interconnect_0:emif_fm_0_emif_usr_clk_clk, rst_controller:clk, tg:emif_usr_clk]
	signal emif_fm_0_pll_ref_clk_out_clk                              : std_logic;                       -- emif_fm_0:pll_ref_clk_out -> local_reset_combiner:clk
	signal emif_cal_emif_calbus_0_calbus_wdata                        : std_logic_vector(31 downto 0);   -- emif_cal:calbus_wdata_0 -> emif_fm_0:calbus_wdata
	signal emif_cal_emif_calbus_0_calbus_address                      : std_logic_vector(19 downto 0);   -- emif_cal:calbus_address_0 -> emif_fm_0:calbus_address
	signal emif_fm_0_emif_calbus_calbus_seq_param_tbl                 : std_logic_vector(4095 downto 0); -- emif_fm_0:calbus_seq_param_tbl -> emif_cal:calbus_seq_param_tbl_0
	signal emif_cal_emif_calbus_0_calbus_read                         : std_logic;                       -- emif_cal:calbus_read_0 -> emif_fm_0:calbus_read
	signal emif_cal_emif_calbus_0_calbus_write                        : std_logic;                       -- emif_cal:calbus_write_0 -> emif_fm_0:calbus_write
	signal emif_fm_0_emif_calbus_calbus_rdata                         : std_logic_vector(31 downto 0);   -- emif_fm_0:calbus_rdata -> emif_cal:calbus_rdata_0
	signal local_reset_source_local_reset_req_local_reset_req         : std_logic;                       -- local_reset_source:local_reset_req -> local_reset_combiner:local_reset_req
	signal local_reset_combiner_local_reset_req_out_0_local_reset_req : std_logic;                       -- local_reset_combiner:local_reset_req_out_0 -> emif_fm_0:local_reset_req
	signal local_reset_combiner_local_reset_status_local_reset_done   : std_logic;                       -- local_reset_combiner:local_reset_done -> local_reset_source:local_reset_done
	signal emif_fm_0_local_reset_status_local_reset_done              : std_logic;                       -- emif_fm_0:local_reset_done -> local_reset_combiner:local_reset_done_in_0
	signal emif_fm_0_mem_mem_reset_n                                  : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_reset_n -> mem:mem_reset_n
	signal emif_fm_0_mem_mem_ba                                       : std_logic_vector(1 downto 0);    -- emif_fm_0:mem_ba -> mem:mem_ba
	signal emif_fm_0_mem_mem_bg                                       : std_logic_vector(1 downto 0);    -- emif_fm_0:mem_bg -> mem:mem_bg
	signal emif_fm_0_mem_mem_ck                                       : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_ck -> mem:mem_ck
	signal emif_fm_0_mem_mem_dqs                                      : std_logic_vector(8 downto 0);    -- [] -> [emif_fm_0:mem_dqs, mem:mem_dqs]
	signal emif_fm_0_mem_mem_act_n                                    : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_act_n -> mem:mem_act_n
	signal emif_fm_0_mem_mem_dq                                       : std_logic_vector(71 downto 0);   -- [] -> [emif_fm_0:mem_dq, mem:mem_dq]
	signal emif_fm_0_mem_mem_cs_n                                     : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_cs_n -> mem:mem_cs_n
	signal emif_fm_0_mem_mem_a                                        : std_logic_vector(16 downto 0);   -- emif_fm_0:mem_a -> mem:mem_a
	signal emif_fm_0_mem_mem_odt                                      : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_odt -> mem:mem_odt
	signal mem_mem_mem_alert_n                                        : std_logic_vector(0 downto 0);    -- mem:mem_alert_n -> emif_fm_0:mem_alert_n
	signal emif_fm_0_mem_mem_dqs_n                                    : std_logic_vector(8 downto 0);    -- [] -> [emif_fm_0:mem_dqs_n, mem:mem_dqs_n]
	signal emif_fm_0_mem_mem_par                                      : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_par -> mem:mem_par
	signal emif_fm_0_mem_mem_dbi_n                                    : std_logic_vector(8 downto 0);    -- [] -> [emif_fm_0:mem_dbi_n, mem:mem_dbi_n]
	signal emif_fm_0_mem_mem_ck_n                                     : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_ck_n -> mem:mem_ck_n
	signal emif_fm_0_mem_mem_cke                                      : std_logic_vector(0 downto 0);    -- emif_fm_0:mem_cke -> mem:mem_cke
	signal emif_fm_0_pll_locked_pll_locked                            : std_logic;                       -- emif_fm_0:pll_locked -> local_reset_combiner:reset_n
	signal emif_fm_0_status_local_cal_fail                            : std_logic;                       -- emif_fm_0:local_cal_fail -> sim_checker:local_cal_fail_0
	signal emif_fm_0_status_local_cal_success                         : std_logic;                       -- emif_fm_0:local_cal_success -> sim_checker:local_cal_success_0
	signal tg_tg_status_0_traffic_gen_fail                            : std_logic;                       -- tg:traffic_gen_fail_0 -> sim_checker:traffic_gen_fail_0
	signal tg_tg_status_0_traffic_gen_timeout                         : std_logic;                       -- tg:traffic_gen_timeout_0 -> sim_checker:traffic_gen_timeout_0
	signal tg_tg_status_0_traffic_gen_pass                            : std_logic;                       -- tg:traffic_gen_pass_0 -> sim_checker:traffic_gen_pass_0
	signal emif_fm_0_emif_usr_reset_n_reset                           : std_logic;                       -- emif_fm_0:emif_usr_reset_n -> [emif_fm_0_emif_usr_reset_n_reset:in, tg:emif_usr_reset_n]
	signal ninit_done_ninit_done_reset                                : std_logic;                       -- ninit_done:ninit_done -> tg:ninit_done
	signal mm_interconnect_0_tg_ctrl_amm_0_waitrequest                : std_logic;                       -- mm_interconnect_0:tg_ctrl_amm_0_waitrequest -> mm_interconnect_0_tg_ctrl_amm_0_waitrequest:in
	signal tg_ctrl_amm_0_readdata                                     : std_logic_vector(575 downto 0);  -- mm_interconnect_0:tg_ctrl_amm_0_readdata -> tg:amm_readdata_0
	signal tg_ctrl_amm_0_read                                         : std_logic;                       -- tg:amm_read_0 -> mm_interconnect_0:tg_ctrl_amm_0_read
	signal tg_ctrl_amm_0_address                                      : std_logic_vector(33 downto 0);   -- tg:amm_address_0 -> mm_interconnect_0:tg_ctrl_amm_0_address
	signal tg_ctrl_amm_0_byteenable                                   : std_logic_vector(71 downto 0);   -- tg:amm_byteenable_0 -> mm_interconnect_0:tg_ctrl_amm_0_byteenable
	signal tg_ctrl_amm_0_readdatavalid                                : std_logic;                       -- mm_interconnect_0:tg_ctrl_amm_0_readdatavalid -> tg:amm_readdatavalid_0
	signal tg_ctrl_amm_0_write                                        : std_logic;                       -- tg:amm_write_0 -> mm_interconnect_0:tg_ctrl_amm_0_write
	signal tg_ctrl_amm_0_writedata                                    : std_logic_vector(575 downto 0);  -- tg:amm_writedata_0 -> mm_interconnect_0:tg_ctrl_amm_0_writedata
	signal tg_ctrl_amm_0_burstcount                                   : std_logic_vector(6 downto 0);    -- tg:amm_burstcount_0 -> mm_interconnect_0:tg_ctrl_amm_0_burstcount
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_readdata            : std_logic_vector(575 downto 0);  -- emif_fm_0:amm_readdata_0 -> mm_interconnect_0:emif_fm_0_ctrl_amm_0_readdata
	signal emif_fm_0_ctrl_amm_0_waitrequest                           : std_logic;                       -- emif_fm_0:amm_ready_0 -> emif_fm_0_ctrl_amm_0_waitrequest:in
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_address             : std_logic_vector(26 downto 0);   -- mm_interconnect_0:emif_fm_0_ctrl_amm_0_address -> emif_fm_0:amm_address_0
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_read                : std_logic;                       -- mm_interconnect_0:emif_fm_0_ctrl_amm_0_read -> emif_fm_0:amm_read_0
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_byteenable          : std_logic_vector(71 downto 0);   -- mm_interconnect_0:emif_fm_0_ctrl_amm_0_byteenable -> emif_fm_0:amm_byteenable_0
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_readdatavalid       : std_logic;                       -- emif_fm_0:amm_readdatavalid_0 -> mm_interconnect_0:emif_fm_0_ctrl_amm_0_readdatavalid
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_write               : std_logic;                       -- mm_interconnect_0:emif_fm_0_ctrl_amm_0_write -> emif_fm_0:amm_write_0
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_writedata           : std_logic_vector(575 downto 0);  -- mm_interconnect_0:emif_fm_0_ctrl_amm_0_writedata -> emif_fm_0:amm_writedata_0
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_burstcount          : std_logic_vector(6 downto 0);    -- mm_interconnect_0:emif_fm_0_ctrl_amm_0_burstcount -> emif_fm_0:amm_burstcount_0
	signal rst_controller_reset_out_reset                             : std_logic;                       -- rst_controller:reset_out -> mm_interconnect_0:tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset
	signal emif_fm_0_emif_usr_reset_n_reset_ports_inv                 : std_logic;                       -- emif_fm_0_emif_usr_reset_n_reset:inv -> rst_controller:reset_in0
	signal tg_ctrl_amm_0_inv                                          : std_logic;                       -- mm_interconnect_0_tg_ctrl_amm_0_waitrequest:inv -> tg:amm_ready_0
	signal mm_interconnect_0_emif_fm_0_ctrl_amm_0_inv                 : std_logic;                       -- emif_fm_0_ctrl_amm_0_waitrequest:inv -> mm_interconnect_0:emif_fm_0_ctrl_amm_0_waitrequest

	for emif_cal : ed_sim_emif_cal_cmp
		use entity ed_sim_emif_cal.ed_sim_emif_cal;
	for emif_fm_0 : ed_sim_emif_fm_0_cmp
		use entity ed_sim_emif_fm_0.ed_sim_emif_fm_0;
	for local_reset_combiner : ed_sim_local_reset_combiner_cmp
		use entity ed_sim_local_reset_combiner.ed_sim_local_reset_combiner;
	for local_reset_source : ed_sim_local_reset_source_cmp
		use entity ed_sim_local_reset_source.ed_sim_local_reset_source;
	for mem : ed_sim_mem_cmp
		use entity ed_sim_mem.ed_sim_mem;
	for ninit_done : ed_sim_ninit_done_cmp
		use entity ed_sim_ninit_done.ed_sim_ninit_done;
	for pll_ref_clk_source : ed_sim_pll_ref_clk_source_cmp
		use entity ed_sim_pll_ref_clk_source.ed_sim_pll_ref_clk_source;
	for sim_checker : ed_sim_sim_checker_cmp
		use entity ed_sim_sim_checker.ed_sim_sim_checker;
	for tg : ed_sim_tg_cmp
		use entity ed_sim_tg.ed_sim_tg;
	for mm_interconnect_0 : ed_sim_altera_mm_interconnect_1920_2l4tnfq_cmp
		use entity altera_mm_interconnect_1920.ed_sim_altera_mm_interconnect_1920_2l4tnfq;
	for rst_controller : altera_reset_controller_cmp
		use entity altera_reset_controller_1921.altera_reset_controller;
begin

	emif_cal : component ed_sim_emif_cal_cmp
		port map (
			calbus_read_0          => emif_cal_emif_calbus_0_calbus_read,         --   emif_calbus_0.calbus_read
			calbus_write_0         => emif_cal_emif_calbus_0_calbus_write,        --                .calbus_write
			calbus_address_0       => emif_cal_emif_calbus_0_calbus_address,      --                .calbus_address
			calbus_wdata_0         => emif_cal_emif_calbus_0_calbus_wdata,        --                .calbus_wdata
			calbus_rdata_0         => emif_fm_0_emif_calbus_calbus_rdata,         --                .calbus_rdata
			calbus_seq_param_tbl_0 => emif_fm_0_emif_calbus_calbus_seq_param_tbl, --                .calbus_seq_param_tbl
			calbus_clk             => emif_cal_emif_calbus_clk_clk                -- emif_calbus_clk.clk
		);

	emif_fm_0 : component ed_sim_emif_fm_0_cmp
		port map (
			local_reset_req      => local_reset_combiner_local_reset_req_out_0_local_reset_req, --    local_reset_req.local_reset_req
			local_reset_done     => emif_fm_0_local_reset_status_local_reset_done,              -- local_reset_status.local_reset_done
			pll_ref_clk          => pll_ref_clk_source_clk_clk,                                 --        pll_ref_clk.clk
			pll_ref_clk_out      => emif_fm_0_pll_ref_clk_out_clk,                              --    pll_ref_clk_out.clk
			pll_locked           => emif_fm_0_pll_locked_pll_locked,                            --         pll_locked.pll_locked
			oct_rzqin            => open,                                                       --                oct.oct_rzqin
			mem_ck               => emif_fm_0_mem_mem_ck,                                       --                mem.mem_ck
			mem_ck_n             => emif_fm_0_mem_mem_ck_n,                                     --                   .mem_ck_n
			mem_a                => emif_fm_0_mem_mem_a,                                        --                   .mem_a
			mem_act_n            => emif_fm_0_mem_mem_act_n,                                    --                   .mem_act_n
			mem_ba               => emif_fm_0_mem_mem_ba,                                       --                   .mem_ba
			mem_bg               => emif_fm_0_mem_mem_bg,                                       --                   .mem_bg
			mem_cke              => emif_fm_0_mem_mem_cke,                                      --                   .mem_cke
			mem_cs_n             => emif_fm_0_mem_mem_cs_n,                                     --                   .mem_cs_n
			mem_odt              => emif_fm_0_mem_mem_odt,                                      --                   .mem_odt
			mem_reset_n          => emif_fm_0_mem_mem_reset_n,                                  --                   .mem_reset_n
			mem_par              => emif_fm_0_mem_mem_par,                                      --                   .mem_par
			mem_alert_n          => mem_mem_mem_alert_n,                                        --                   .mem_alert_n
			mem_dqs              => emif_fm_0_mem_mem_dqs,                                      --                   .mem_dqs
			mem_dqs_n            => emif_fm_0_mem_mem_dqs_n,                                    --                   .mem_dqs_n
			mem_dq               => emif_fm_0_mem_mem_dq,                                       --                   .mem_dq
			mem_dbi_n            => emif_fm_0_mem_mem_dbi_n,                                    --                   .mem_dbi_n
			local_cal_success    => emif_fm_0_status_local_cal_success,                         --             status.local_cal_success
			local_cal_fail       => emif_fm_0_status_local_cal_fail,                            --                   .local_cal_fail
			emif_usr_reset_n     => emif_fm_0_emif_usr_reset_n_reset,                           --   emif_usr_reset_n.reset_n
			emif_usr_clk         => emif_fm_0_emif_usr_clk_clk,                                 --       emif_usr_clk.clk
			amm_ready_0          => emif_fm_0_ctrl_amm_0_waitrequest,                           --         ctrl_amm_0.waitrequest_n
			amm_read_0           => mm_interconnect_0_emif_fm_0_ctrl_amm_0_read,                --                   .read
			amm_write_0          => mm_interconnect_0_emif_fm_0_ctrl_amm_0_write,               --                   .write
			amm_address_0        => mm_interconnect_0_emif_fm_0_ctrl_amm_0_address,             --                   .address
			amm_readdata_0       => mm_interconnect_0_emif_fm_0_ctrl_amm_0_readdata,            --                   .readdata
			amm_writedata_0      => mm_interconnect_0_emif_fm_0_ctrl_amm_0_writedata,           --                   .writedata
			amm_burstcount_0     => mm_interconnect_0_emif_fm_0_ctrl_amm_0_burstcount,          --                   .burstcount
			amm_byteenable_0     => mm_interconnect_0_emif_fm_0_ctrl_amm_0_byteenable,          --                   .byteenable
			amm_readdatavalid_0  => mm_interconnect_0_emif_fm_0_ctrl_amm_0_readdatavalid,       --                   .readdatavalid
			calbus_read          => emif_cal_emif_calbus_0_calbus_read,                         --        emif_calbus.calbus_read
			calbus_write         => emif_cal_emif_calbus_0_calbus_write,                        --                   .calbus_write
			calbus_address       => emif_cal_emif_calbus_0_calbus_address,                      --                   .calbus_address
			calbus_wdata         => emif_cal_emif_calbus_0_calbus_wdata,                        --                   .calbus_wdata
			calbus_rdata         => emif_fm_0_emif_calbus_calbus_rdata,                         --                   .calbus_rdata
			calbus_seq_param_tbl => emif_fm_0_emif_calbus_calbus_seq_param_tbl,                 --                   .calbus_seq_param_tbl
			calbus_clk           => emif_cal_emif_calbus_clk_clk                                --    emif_calbus_clk.clk
		);

	local_reset_combiner : component ed_sim_local_reset_combiner_cmp
		port map (
			local_reset_req_out_0 => local_reset_combiner_local_reset_req_out_0_local_reset_req, --   local_reset_req_out_0.local_reset_req
			local_reset_done_in_0 => emif_fm_0_local_reset_status_local_reset_done,              -- local_reset_status_in_0.local_reset_done
			clk                   => emif_fm_0_pll_ref_clk_out_clk,                              --             generic_clk.clk
			reset_n               => emif_fm_0_pll_locked_pll_locked,                            -- generic_conduit_reset_n.pll_locked
			local_reset_req       => local_reset_source_local_reset_req_local_reset_req,         --         local_reset_req.local_reset_req
			local_reset_done      => local_reset_combiner_local_reset_status_local_reset_done    --      local_reset_status.local_reset_done
		);

	local_reset_source : component ed_sim_local_reset_source_cmp
		port map (
			local_reset_req  => local_reset_source_local_reset_req_local_reset_req,       --    local_reset_req.local_reset_req
			local_reset_done => local_reset_combiner_local_reset_status_local_reset_done  -- local_reset_status.local_reset_done
		);

	mem : component ed_sim_mem_cmp
		port map (
			mem_ck      => emif_fm_0_mem_mem_ck,      -- mem.mem_ck
			mem_ck_n    => emif_fm_0_mem_mem_ck_n,    --    .mem_ck_n
			mem_a       => emif_fm_0_mem_mem_a,       --    .mem_a
			mem_act_n   => emif_fm_0_mem_mem_act_n,   --    .mem_act_n
			mem_ba      => emif_fm_0_mem_mem_ba,      --    .mem_ba
			mem_bg      => emif_fm_0_mem_mem_bg,      --    .mem_bg
			mem_cke     => emif_fm_0_mem_mem_cke,     --    .mem_cke
			mem_cs_n    => emif_fm_0_mem_mem_cs_n,    --    .mem_cs_n
			mem_odt     => emif_fm_0_mem_mem_odt,     --    .mem_odt
			mem_reset_n => emif_fm_0_mem_mem_reset_n, --    .mem_reset_n
			mem_par     => emif_fm_0_mem_mem_par,     --    .mem_par
			mem_alert_n => mem_mem_mem_alert_n,       --    .mem_alert_n
			mem_dqs     => emif_fm_0_mem_mem_dqs,     --    .mem_dqs
			mem_dqs_n   => emif_fm_0_mem_mem_dqs_n,   --    .mem_dqs_n
			mem_dq      => emif_fm_0_mem_mem_dq,      --    .mem_dq
			mem_dbi_n   => emif_fm_0_mem_mem_dbi_n    --    .mem_dbi_n
		);

	ninit_done : component ed_sim_ninit_done_cmp
		port map (
			ninit_done => ninit_done_ninit_done_reset  -- ninit_done.reset
		);

	pll_ref_clk_source : component ed_sim_pll_ref_clk_source_cmp
		port map (
			clk => pll_ref_clk_source_clk_clk  -- clk.clk
		);

	sim_checker : component ed_sim_sim_checker_cmp
		port map (
			traffic_gen_pass_0    => tg_tg_status_0_traffic_gen_pass,      -- tg_status_0.traffic_gen_pass
			traffic_gen_fail_0    => tg_tg_status_0_traffic_gen_fail,      --            .traffic_gen_fail
			traffic_gen_timeout_0 => tg_tg_status_0_traffic_gen_timeout,   --            .traffic_gen_timeout
			traffic_gen_pass      => sim_checker_traffic_gen_pass,         --   tg_status.traffic_gen_pass
			traffic_gen_fail      => sim_checker_traffic_gen_fail,         --            .traffic_gen_fail
			traffic_gen_timeout   => sim_checker_traffic_gen_timeout,      --            .traffic_gen_timeout
			local_cal_success_0   => emif_fm_0_status_local_cal_success,   --    status_0.local_cal_success
			local_cal_fail_0      => emif_fm_0_status_local_cal_fail,      --            .local_cal_fail
			local_cal_success     => cal_status_checker_local_cal_success, --      status.local_cal_success
			local_cal_fail        => cal_status_checker_local_cal_fail     --            .local_cal_fail
		);

	tg : component ed_sim_tg_cmp
		port map (
			emif_usr_reset_n      => emif_fm_0_emif_usr_reset_n_reset,   -- emif_usr_reset_n.reset_n
			ninit_done            => ninit_done_ninit_done_reset,        --       ninit_done.reset
			emif_usr_clk          => emif_fm_0_emif_usr_clk_clk,         --     emif_usr_clk.clk
			amm_ready_0           => tg_ctrl_amm_0_inv,                  --       ctrl_amm_0.waitrequest_n
			amm_read_0            => tg_ctrl_amm_0_read,                 --                 .read
			amm_write_0           => tg_ctrl_amm_0_write,                --                 .write
			amm_address_0         => tg_ctrl_amm_0_address,              --                 .address
			amm_readdata_0        => tg_ctrl_amm_0_readdata,             --                 .readdata
			amm_writedata_0       => tg_ctrl_amm_0_writedata,            --                 .writedata
			amm_burstcount_0      => tg_ctrl_amm_0_burstcount,           --                 .burstcount
			amm_byteenable_0      => tg_ctrl_amm_0_byteenable,           --                 .byteenable
			amm_readdatavalid_0   => tg_ctrl_amm_0_readdatavalid,        --                 .readdatavalid
			traffic_gen_pass_0    => tg_tg_status_0_traffic_gen_pass,    --      tg_status_0.traffic_gen_pass
			traffic_gen_fail_0    => tg_tg_status_0_traffic_gen_fail,    --                 .traffic_gen_fail
			traffic_gen_timeout_0 => tg_tg_status_0_traffic_gen_timeout  --                 .traffic_gen_timeout
		);

	mm_interconnect_0 : component ed_sim_altera_mm_interconnect_1920_2l4tnfq_cmp
		port map (
			tg_ctrl_amm_0_address                                      => tg_ctrl_amm_0_address,                                --                                        tg_ctrl_amm_0.address
			tg_ctrl_amm_0_waitrequest                                  => mm_interconnect_0_tg_ctrl_amm_0_waitrequest,          --                                                     .waitrequest
			tg_ctrl_amm_0_burstcount                                   => tg_ctrl_amm_0_burstcount,                             --                                                     .burstcount
			tg_ctrl_amm_0_byteenable                                   => tg_ctrl_amm_0_byteenable,                             --                                                     .byteenable
			tg_ctrl_amm_0_read                                         => tg_ctrl_amm_0_read,                                   --                                                     .read
			tg_ctrl_amm_0_readdata                                     => tg_ctrl_amm_0_readdata,                               --                                                     .readdata
			tg_ctrl_amm_0_readdatavalid                                => tg_ctrl_amm_0_readdatavalid,                          --                                                     .readdatavalid
			tg_ctrl_amm_0_write                                        => tg_ctrl_amm_0_write,                                  --                                                     .write
			tg_ctrl_amm_0_writedata                                    => tg_ctrl_amm_0_writedata,                              --                                                     .writedata
			emif_fm_0_ctrl_amm_0_address                               => mm_interconnect_0_emif_fm_0_ctrl_amm_0_address,       --                                 emif_fm_0_ctrl_amm_0.address
			emif_fm_0_ctrl_amm_0_write                                 => mm_interconnect_0_emif_fm_0_ctrl_amm_0_write,         --                                                     .write
			emif_fm_0_ctrl_amm_0_read                                  => mm_interconnect_0_emif_fm_0_ctrl_amm_0_read,          --                                                     .read
			emif_fm_0_ctrl_amm_0_readdata                              => mm_interconnect_0_emif_fm_0_ctrl_amm_0_readdata,      --                                                     .readdata
			emif_fm_0_ctrl_amm_0_writedata                             => mm_interconnect_0_emif_fm_0_ctrl_amm_0_writedata,     --                                                     .writedata
			emif_fm_0_ctrl_amm_0_burstcount                            => mm_interconnect_0_emif_fm_0_ctrl_amm_0_burstcount,    --                                                     .burstcount
			emif_fm_0_ctrl_amm_0_byteenable                            => mm_interconnect_0_emif_fm_0_ctrl_amm_0_byteenable,    --                                                     .byteenable
			emif_fm_0_ctrl_amm_0_readdatavalid                         => mm_interconnect_0_emif_fm_0_ctrl_amm_0_readdatavalid, --                                                     .readdatavalid
			emif_fm_0_ctrl_amm_0_waitrequest                           => mm_interconnect_0_emif_fm_0_ctrl_amm_0_inv,           --                                                     .waitrequest
			tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset.reset
			emif_fm_0_emif_usr_clk_clk                                 => emif_fm_0_emif_usr_clk_clk                            --                               emif_fm_0_emif_usr_clk.clk
		);

	rst_controller : component altera_reset_controller_cmp
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "both",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => emif_fm_0_emif_usr_reset_n_reset_ports_inv, -- reset_in0.reset
			clk            => emif_fm_0_emif_usr_clk_clk,                 --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_in1      => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	emif_fm_0_emif_usr_reset_n_reset_ports_inv <= not emif_fm_0_emif_usr_reset_n_reset;

	tg_ctrl_amm_0_inv <= not mm_interconnect_0_tg_ctrl_amm_0_waitrequest;

	mm_interconnect_0_emif_fm_0_ctrl_amm_0_inv <= not emif_fm_0_ctrl_amm_0_waitrequest;

end architecture rtl; -- of ed_sim
