-- PCIE_HIP_FDAS_altera_merlin_burst_adapter_altera_avalon_st_pipeline_stage_1922_wyh7ycq.vhd

-- Generated using ACDS version 22.2 94

library IEEE;
library altera_avalon_st_pipeline_stage_1920;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PCIE_HIP_FDAS_altera_merlin_burst_adapter_altera_avalon_st_pipeline_stage_1922_wyh7ycq is
	generic (
		SYMBOLS_PER_BEAT : integer := 1;
		BITS_PER_SYMBOL  : integer := 147;
		USE_PACKETS      : integer := 1;
		USE_EMPTY        : integer := 0;
		EMPTY_WIDTH      : integer := 0;
		CHANNEL_WIDTH    : integer := 1;
		PACKET_WIDTH     : integer := 2;
		ERROR_WIDTH      : integer := 0;
		PIPELINE_READY   : integer := 1;
		SYNC_RESET       : integer := 1
	);
	port (
		clk               : in  std_logic                      := '0';             --       cr0.clk
		reset             : in  std_logic                      := '0';             -- cr0_reset.reset
		in_ready          : out std_logic;                                         --     sink0.ready
		in_valid          : in  std_logic                      := '0';             --          .valid
		in_startofpacket  : in  std_logic                      := '0';             --          .startofpacket
		in_endofpacket    : in  std_logic                      := '0';             --          .endofpacket
		in_data           : in  std_logic_vector(146 downto 0) := (others => '0'); --          .data
		in_channel        : in  std_logic_vector(0 downto 0)   := (others => '0'); --          .channel
		out_ready         : in  std_logic                      := '0';             --   source0.ready
		out_valid         : out std_logic;                                         --          .valid
		out_startofpacket : out std_logic;                                         --          .startofpacket
		out_endofpacket   : out std_logic;                                         --          .endofpacket
		out_data          : out std_logic_vector(146 downto 0);                    --          .data
		out_channel       : out std_logic_vector(0 downto 0)                       --          .channel
	);
end entity PCIE_HIP_FDAS_altera_merlin_burst_adapter_altera_avalon_st_pipeline_stage_1922_wyh7ycq;

architecture rtl of PCIE_HIP_FDAS_altera_merlin_burst_adapter_altera_avalon_st_pipeline_stage_1922_wyh7ycq is
	component PCIE_HIP_FDAS_altera_avalon_st_pipeline_stage_1920_zterisq_cmp is
		generic (
			SYMBOLS_PER_BEAT : integer := 1;
			BITS_PER_SYMBOL  : integer := 8;
			USE_PACKETS      : integer := 0;
			USE_EMPTY        : integer := 0;
			EMPTY_WIDTH      : integer := 0;
			CHANNEL_WIDTH    : integer := 0;
			PACKET_WIDTH     : integer := 0;
			ERROR_WIDTH      : integer := 0;
			PIPELINE_READY   : integer := 1;
			SYNC_RESET       : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_ready          : out std_logic;                                         -- ready
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_data           : in  std_logic_vector(146 downto 0) := (others => 'X'); -- data
			in_channel        : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- channel
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_valid         : out std_logic;                                         -- valid
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_data          : out std_logic_vector(146 downto 0);                    -- data
			out_channel       : out std_logic_vector(0 downto 0);                      -- channel
			in_empty          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- empty
			out_empty         : out std_logic_vector(0 downto 0);                      -- empty
			out_error         : out std_logic_vector(0 downto 0);                      -- error
			in_error          : in  std_logic_vector(0 downto 0)   := (others => 'X')  -- error
		);
	end component PCIE_HIP_FDAS_altera_avalon_st_pipeline_stage_1920_zterisq_cmp;

	for my_altera_avalon_st_pipeline_stage : PCIE_HIP_FDAS_altera_avalon_st_pipeline_stage_1920_zterisq_cmp
		use entity altera_avalon_st_pipeline_stage_1920.PCIE_HIP_FDAS_altera_avalon_st_pipeline_stage_1920_zterisq;
begin

	my_altera_avalon_st_pipeline_stage : component PCIE_HIP_FDAS_altera_avalon_st_pipeline_stage_1920_zterisq_cmp
		generic map (
			SYMBOLS_PER_BEAT => SYMBOLS_PER_BEAT,
			BITS_PER_SYMBOL  => BITS_PER_SYMBOL,
			USE_PACKETS      => USE_PACKETS,
			USE_EMPTY        => USE_EMPTY,
			EMPTY_WIDTH      => EMPTY_WIDTH,
			CHANNEL_WIDTH    => CHANNEL_WIDTH,
			PACKET_WIDTH     => PACKET_WIDTH,
			ERROR_WIDTH      => ERROR_WIDTH,
			PIPELINE_READY   => PIPELINE_READY,
			SYNC_RESET       => SYNC_RESET
		)
		port map (
			clk               => clk,               --       cr0.clk
			reset             => reset,             -- cr0_reset.reset
			in_ready          => in_ready,          --     sink0.ready
			in_valid          => in_valid,          --          .valid
			in_startofpacket  => in_startofpacket,  --          .startofpacket
			in_endofpacket    => in_endofpacket,    --          .endofpacket
			in_data           => in_data,           --          .data
			in_channel        => in_channel,        --          .channel
			out_ready         => out_ready,         --   source0.ready
			out_valid         => out_valid,         --          .valid
			out_startofpacket => out_startofpacket, --          .startofpacket
			out_endofpacket   => out_endofpacket,   --          .endofpacket
			out_data          => out_data,          --          .data
			out_channel       => out_channel,       --          .channel
			in_empty          => "0",               -- (terminated)
			out_empty         => open,              -- (terminated)
			out_error         => open,              -- (terminated)
			in_error          => "0"                -- (terminated)
		);

end architecture rtl; -- of PCIE_HIP_FDAS_altera_merlin_burst_adapter_altera_avalon_st_pipeline_stage_1922_wyh7ycq
