----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.conv_fft_str.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 18:56:38 11/07/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library conv_lib;

entity conv_fft_str is
  generic( 
    dbits_g     : natural;
    depth_g     : natural;
    abits_g     : natural;
    pages_g     : natural;    -- lte 2**pgbits_g
    pgbits_g    : natural;
    loop_g      : natural;    -- number of output frame repeats lte 2**loop_bits_g 
    loop_bits_g : natural
  );
  port( 
    CLK_SYS        : in     std_logic;
    RST_SYS_N      : in     std_logic;
    RDATAOUT       : out    std_logic_vector (dbits_g-1 downto 0);
    IDATAOUT       : out    std_logic_vector (dbits_g-1 downto 0);
    VALIDOUT       : out    std_logic;
    SOFOUT         : out    std_logic;
    EOFOUT         : out    std_logic;
    LOOP_ADDROUT   : out    std_logic_vector (loop_bits_g-1 downto 0);
    READYOUT       : out    std_logic;
    COEF_RDENOUT   : out    std_logic_vector (loop_g-1 downto 0);
    COEF_RDADDROUT : out    std_logic_vector (abits_g-1 downto 0);
    RDATA          : in     std_logic_vector (dbits_g-1 downto 0);
    IDATA          : in     std_logic_vector (dbits_g-1 downto 0);
    VALID          : in     std_logic;
    SOF            : in     std_logic;
    EOF            : in     std_logic;
    LOOP_NUM       : in     std_logic_vector (loop_bits_g downto 0);
    CONV_ENABLE    : in     std_logic;
    SYNC           : in     std_logic;
    READY          : in     std_logic_vector (loop_g-1 downto 0);
    CLK_MC         : in     std_logic;
    RST_MC_N       : in     std_logic;
    MCADDR         : in     std_logic_vector (abits_g downto 0);
    MCRDEN         : in     std_logic;
    MCDATAOUT      : out    std_logic_vector (dbits_g-1 downto 0);
    DONEOUT        : out    std_logic;
    OVERFLOW       : out    std_logic
  );

-- Declarations

end entity conv_fft_str ;

