----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity ctrl_lib.ctrl.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 11:59:37 17/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ctrl is
  port( 
    cld_done       : in     std_logic;
    clk_mc         : in     std_logic;
    clk_sys        : in     std_logic;
    conv_done      : in     std_logic;
    conv_fft_ready : in     std_logic;
    conv_waitreq   : in     std_logic;
    conv_wr_en     : in     std_logic;
    hsum_done      : in     std_logic;
    hsum_rd_en     : in     std_logic;
    hsum_valid     : in     std_logic;
    hsum_waitreq   : in     std_logic;
    mcaddr         : in     std_logic_vector (18 downto 0);
    mcdatain       : in     std_logic_vector (31 downto 0);
    mcms           : in     std_logic;
    mcrwn          : in     std_logic;
    rst_mc_n       : in     std_logic;
    rst_sys_n      : in     std_logic;
    cld_enable     : out    std_logic;
    cld_page       : out    std_logic_vector (31 downto 0);
    cld_trigger    : out    std_logic;
    conv_enable    : out    std_logic;
    conv_page      : out    std_logic_vector (31 downto 0);
    conv_trigger   : out    std_logic;
    fop_sample_num : out    std_logic_vector (22 downto 0);
    hsum_enable    : out    std_logic;
    hsum_page      : out    std_logic_vector (31 downto 0);
    hsum_trigger   : out    std_logic;
    ifft_loop_num  : out    std_logic_vector (5 downto 0);
    mcdataout      : out    std_logic_vector (31 downto 0);
    overlap_size   : out    std_logic_vector (9 downto 0)
  );

-- Declarations

end entity ctrl ;

