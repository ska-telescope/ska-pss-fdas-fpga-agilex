----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity pcif_lib.pcif.symbol
--
-- Created:
--          by - droogm.UNKNOWN (COVNETICSDT7)
--          at - 11:57:51 03/11/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY pcif IS
   PORT( 
      clk_mc                   : IN     std_logic;
      clk_pcie                 : IN     std_logic;
      mcdataout                : IN     std_logic_vector (31 DOWNTO 0);
      rst_mc_n                 : IN     std_logic;
      rst_pcie_n               : IN     std_logic;
      rxm_address              : IN     std_logic_vector (21 DOWNTO 0);
      rxm_byte_enable          : IN     std_logic_vector (3 DOWNTO 0);
      rxm_read                 : IN     std_logic;
      rxm_write                : IN     std_logic;
      rxm_write_data           : IN     std_logic_vector (31 DOWNTO 0);
      mcaddr                   : OUT    std_logic_vector (21 DOWNTO 0);
      mccs                     : OUT    std_logic;
      mcdatain                 : OUT    std_logic_vector (31 DOWNTO 0);
      mcrwn                    : OUT    std_logic;
      rxm_read_data            : OUT    std_logic_vector (31 DOWNTO 0);
      rxm_read_data_vald       : OUT    std_logic;
      rxm_response             : OUT    std_logic_vector (1 DOWNTO 0);
      rxm_wait_request         : OUT    std_logic;
      rxm_write_response_valid : OUT    std_logic
   );

-- Declarations

END pcif ;

