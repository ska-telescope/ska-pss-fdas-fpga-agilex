----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2022 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.conv_mult.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT11)
--          at - 14:09:22 22/04/2022
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.2a (Build 3)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity conv_mult is
  port( 
    CLK_SYS      : in     std_logic;
    ICOEF        : in     std_logic_vector (31 downto 0);
    ICOEFCONJ    : in     std_logic_vector (31 downto 0);
    IDATA        : in     std_logic_vector (31 downto 0);
    RCOEF        : in     std_logic_vector (31 downto 0);
    RCOEFCONJ    : in     std_logic_vector (31 downto 0);
    RDATA        : in     std_logic_vector (31 downto 0);
    RST_SYS_N    : in     std_logic;
    VALID        : in     std_logic;
    IDATACONJOUT : out    std_logic_vector (31 downto 0);  -- result
    IDATAOUT     : out    std_logic_vector (31 downto 0);
    RDATACONJOUT : out    std_logic_vector (31 downto 0);  -- result
    RDATAOUT     : out    std_logic_vector (31 downto 0)
  );

-- Declarations

end entity conv_mult ;

