----------------------------------------------------------------------------
--       __
--    ,/'__`\                             _     _
--   ,/ /  )_)   _   _   _   ___     __  | |__ (_)   __    ___
--   ( (    _  /' `\\ \ / //' _ `\ /'__`\|  __)| | /'__`)/',__)
--   '\ \__) )( (_) )\ ' / | ( ) |(  ___/| |_, | |( (___ \__, \
--    '\___,/  \___/  \_/  (_) (_)`\____)(___,)(_)`\___,)(____/
--
-- Copyright (c) Covnetics Limited 2017 All Rights Reserved. The information
-- contained herein remains the property of Covnetics Limited and may not be
-- copied or reproduced in any format or medium without the written consent
-- of Covnetics Limited.
--
----------------------------------------------------------------------------
-- VHDL Entity conv_lib.retime.symbol
--
-- Created:
--          by - taylorj.UNKNOWN (COVNETICSDT1)
--          at - 10:22:09 12/06/2017
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity retime is
  generic( 
    dataw_g  : natural;
    stages_g : natural
  );
  port( 
    DATA    : in     std_logic_vector (dataw_g-1 downto 0);
    DE      : in     std_logic;
    SYNC    : in     std_logic;
    CLK     : in     std_logic;
    CLKEN   : in     std_logic;
    RST_N   : in     std_logic;
    DATAOUT : out    std_logic_vector (dataw_g-1 downto 0);
    DEOUT   : out    std_logic
  );

-- Declarations

end entity retime ;
